library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn7411_tb is
end sn7411_tb;

architecture testbench of sn7411_tb is

begin

--  uut : sn7411 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
