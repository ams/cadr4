library ieee;
use ieee.std_logic_1164.all;

entity cadr_vma is
  port (
    \-srcvma\       : in     std_logic;
    \-vmaenb\       : in     std_logic;
    \-vmas0\        : in     std_logic;
    \-vmas10\       : in     std_logic;
    \-vmas11\       : in     std_logic;
    \-vmas12\       : in     std_logic;
    \-vmas13\       : in     std_logic;
    \-vmas14\       : in     std_logic;
    \-vmas15\       : in     std_logic;
    \-vmas16\       : in     std_logic;
    \-vmas17\       : in     std_logic;
    \-vmas18\       : in     std_logic;
    \-vmas19\       : in     std_logic;
    \-vmas1\        : in     std_logic;
    \-vmas20\       : in     std_logic;
    \-vmas21\       : in     std_logic;
    \-vmas22\       : in     std_logic;
    \-vmas23\       : in     std_logic;
    \-vmas24\       : in     std_logic;
    \-vmas25\       : in     std_logic;
    \-vmas26\       : in     std_logic;
    \-vmas27\       : in     std_logic;
    \-vmas28\       : in     std_logic;
    \-vmas29\       : in     std_logic;
    \-vmas2\        : in     std_logic;
    \-vmas30\       : in     std_logic;
    \-vmas31\       : in     std_logic;
    \-vmas3\        : in     std_logic;
    \-vmas4\        : in     std_logic;
    \-vmas5\        : in     std_logic;
    \-vmas6\        : in     std_logic;
    \-vmas7\        : in     std_logic;
    \-vmas8\        : in     std_logic;
    \-vmas9\        : in     std_logic;
    clk1a           : in     std_logic;
    clk2a           : in     std_logic;
    clk2c           : in     std_logic;
    tse2            : in     std_logic;
    \-vma0\         : out    std_logic;
    \-vma10\        : out    std_logic;
    \-vma11\        : out    std_logic;
    \-vma12\        : out    std_logic;
    \-vma13\        : out    std_logic;
    \-vma14\        : out    std_logic;
    \-vma15\        : out    std_logic;
    \-vma16\        : out    std_logic;
    \-vma17\        : out    std_logic;
    \-vma18\        : out    std_logic;
    \-vma19\        : out    std_logic;
    \-vma1\         : out    std_logic;
    \-vma20\        : out    std_logic;
    \-vma21\        : out    std_logic;
    \-vma22\        : out    std_logic;
    \-vma23\        : out    std_logic;
    \-vma24\        : out    std_logic;
    \-vma25\        : out    std_logic;
    \-vma26\        : out    std_logic;
    \-vma27\        : out    std_logic;
    \-vma28\        : out    std_logic;
    \-vma29\        : out    std_logic;
    \-vma2\         : out    std_logic;
    \-vma30\        : out    std_logic;
    \-vma31\        : out    std_logic;
    \-vma3\         : out    std_logic;
    \-vma4\         : out    std_logic;
    \-vma5\         : out    std_logic;
    \-vma6\         : out    std_logic;
    \-vma7\         : out    std_logic;
    \-vma8\         : out    std_logic;
    \-vma9\         : out    std_logic;
    \-vmadrive\     : out    std_logic;
    mf0             : out    std_logic;
    mf1             : out    std_logic;
    mf10            : out    std_logic;
    mf11            : out    std_logic;
    mf12            : out    std_logic;
    mf13            : out    std_logic;
    mf14            : out    std_logic;
    mf15            : out    std_logic;
    mf16            : out    std_logic;
    mf17            : out    std_logic;
    mf18            : out    std_logic;
    mf19            : out    std_logic;
    mf2             : out    std_logic;
    mf20            : out    std_logic;
    mf21            : out    std_logic;
    mf22            : out    std_logic;
    mf23            : out    std_logic;
    mf24            : out    std_logic;
    mf25            : out    std_logic;
    mf26            : out    std_logic;
    mf27            : out    std_logic;
    mf28            : out    std_logic;
    mf29            : out    std_logic;
    mf3             : out    std_logic;
    mf30            : out    std_logic;
    mf31            : out    std_logic;
    mf4             : out    std_logic;
    mf5             : out    std_logic;
    mf6             : out    std_logic;
    mf7             : out    std_logic;
    mf8             : out    std_logic;
    mf9             : out    std_logic;
    srcvma          : out    std_logic
  );
end entity;
