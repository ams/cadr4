library ieee;
use ieee.std_logic_1164.all;

entity cadr1_uba is
  port (
    \-ub adr0\      : in     std_logic;
    \-ub adr10\     : in     std_logic;
    \-ub adr11\     : in     std_logic;
    \-ub adr12\     : in     std_logic;
    \-ub adr13\     : in     std_logic;
    \-ub adr14\     : in     std_logic;
    \-ub adr15\     : in     std_logic;
    \-ub adr16\     : in     std_logic;
    \-ub adr17\     : in     std_logic;
    \-ub adr1\      : in     std_logic;
    \-ub adr2\      : in     std_logic;
    \-ub adr3\      : in     std_logic;
    \-ub adr4\      : in     std_logic;
    \-ub adr5\      : in     std_logic;
    \-ub adr6\      : in     std_logic;
    \-ub adr7\      : in     std_logic;
    \-ub adr8\      : in     std_logic;
    \-ub adr9\      : in     std_logic;
    \-ub c1\        : in     std_logic;
    \-ubadrive\     : in     std_logic;
    \c1 in\         : in     std_logic;
    \c1 out\        : in     std_logic;
    uao1            : in     std_logic;
    uao10           : in     std_logic;
    uao11           : in     std_logic;
    uao12           : in     std_logic;
    uao13           : in     std_logic;
    uao14           : in     std_logic;
    uao15           : in     std_logic;
    uao16           : in     std_logic;
    uao17           : in     std_logic;
    uao2            : in     std_logic;
    uao3            : in     std_logic;
    uao4            : in     std_logic;
    uao5            : in     std_logic;
    uao6            : in     std_logic;
    uao7            : in     std_logic;
    uao8            : in     std_logic;
    uao9            : in     std_logic;
    uba0            : in     std_logic;
    uba1            : in     std_logic;
    uba10           : in     std_logic;
    uba11           : in     std_logic;
    uba12           : in     std_logic;
    uba13           : in     std_logic;
    uba14           : in     std_logic;
    uba15           : in     std_logic;
    uba16           : in     std_logic;
    uba17           : in     std_logic;
    uba2            : in     std_logic;
    uba3            : in     std_logic;
    uba4            : in     std_logic;
    uba5            : in     std_logic;
    uba6            : in     std_logic;
    uba7            : in     std_logic;
    uba8            : in     std_logic;
    uba9            : in     std_logic;
    \-uba 12\       : out    std_logic;
    \-uba 14\       : out    std_logic;
    \-uba 15\       : out    std_logic;
    \-uba 7\        : out    std_logic;
    \-uba 8\        : out    std_logic;
    \-uba 9\        : out    std_logic
  );
end entity cadr1_uba;
