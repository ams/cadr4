library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sip220_330_8 is
  port (
    r2 : out std_logic;
    r3 : out std_logic;
    r4 : out std_logic;
    r5 : out std_logic;
    r6 : out std_logic;
    r7 : out std_logic
    );
end;

architecture ttl of sip220_330_8 is
begin
  r2 <= '1'; r3 <= '1'; r4 <= '1';
  r5 <= '1'; r6 <= '1'; r7 <= '1';
end;
