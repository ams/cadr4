library ieee;
use ieee.std_logic_1164.all;

entity vmemdr is
  port (
    \-mapdrive\ : out std_logic;
    \-pfw\      : in  std_logic;
    mf24        : out std_logic;
    \-pfr\      : in  std_logic;
    mf25        : out std_logic;
    hi12        : in  std_logic;
    mf26        : out std_logic;
    \-vmap4\    : in  std_logic;
    mf27        : out std_logic;
    \-vmap3\    : in  std_logic;
    mf28        : out std_logic;
    \-vmap2\    : in  std_logic;
    mf29        : out std_logic;
    \-vmap1\    : in  std_logic;
    mf30        : out std_logic;
    \-vmap0\    : in  std_logic;
    mf31        : out std_logic;
    \-vmo15\    : in  std_logic;
    mf8         : out std_logic;
    \-vmo14\    : in  std_logic;
    mf9         : out std_logic;
    \-vmo13\    : in  std_logic;
    mf10        : out std_logic;
    \-vmo12\    : in  std_logic;
    mf11        : out std_logic;
    \-vmo11\    : in  std_logic;
    mf12        : out std_logic;
    \-vmo10\    : in  std_logic;
    mf13        : out std_logic;
    \-vmo9\     : in  std_logic;
    mf14        : out std_logic;
    \-vmo8\     : in  std_logic;
    mf15        : out std_logic;
    \-vmo23\    : in  std_logic;
    mf16        : out std_logic;
    \-vmo22\    : in  std_logic;
    mf17        : out std_logic;
    \-vmo21\    : in  std_logic;
    mf18        : out std_logic;
    \-vmo20\    : in  std_logic;
    mf19        : out std_logic;
    \-vmo19\    : in  std_logic;
    mf20        : out std_logic;
    \-vmo18\    : in  std_logic;
    mf21        : out std_logic;
    \-vmo17\    : in  std_logic;
    mf22        : out std_logic;
    \-vmo16\    : in  std_logic;
    mf23        : out std_logic;
    tse1a       : in  std_logic;
    srcmap      : out std_logic;
    \-vmo7\     : in  std_logic;
    mf0         : out std_logic;
    \-vmo6\     : in  std_logic;
    mf1         : out std_logic;
    \-vmo5\     : in  std_logic;
    mf2         : out std_logic;
    \-vmo4\     : in  std_logic;
    mf3         : out std_logic;
    \-vmo3\     : in  std_logic;
    mf4         : out std_logic;
    \-vmo2\     : in  std_logic;
    mf5         : out std_logic;
    \-vmo1\     : in  std_logic;
    mf6         : out std_logic;
    \-vmo0\     : in  std_logic;
    mf7         : out std_logic;
    gnd         : in  std_logic;
    \-lvmo23\   : out std_logic;
    \-lvmo22\   : out std_logic;
    \-pma21\    : out std_logic;
    \-pma20\    : out std_logic;
    memstart    : in  std_logic;
    \-pma19\    : out std_logic;
    \-pma18\    : out std_logic;
    \-pma17\    : out std_logic;
    \-pma16\    : out std_logic;
    \-pma15\    : out std_logic;
    \-pma14\    : out std_logic;
    \-pma13\    : out std_logic;
    \-pma12\    : out std_logic;
    \-pma11\    : out std_logic;
    \-pma10\    : out std_logic;
    \-pma9\     : out std_logic;
    \-pma8\     : out std_logic;
    \-vma6\     : in  std_logic;
    \-vma5\     : in  std_logic;
    \-vma4\     : in  std_logic;
    \-vma3\     : in  std_logic;
    \-vma2\     : in  std_logic;
    \-vma1\     : in  std_logic;
    \-vma0\     : in  std_logic;
    \-vma7\     : in  std_logic;
    \-adrpar\   : out std_logic;
    \-srcmap\   : in  std_logic);
end;
