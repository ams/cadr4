library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_md is
  port (
    \-mddrive\  : out std_logic;
    \-md31\     : out std_logic;
    mf24        : out std_logic;
    \-md30\     : out std_logic;
    mf25        : out std_logic;
    \-md29\     : out std_logic;
    mf26        : out std_logic;
    \-md28\     : out std_logic;
    mf27        : out std_logic;
    \-md27\     : out std_logic;
    mf28        : out std_logic;
    \-md26\     : out std_logic;
    mf29        : out std_logic;
    \-md25\     : out std_logic;
    mf30        : out std_logic;
    \-md24\     : out std_logic;
    mf31        : out std_logic;
    \-md23\     : out std_logic;
    mf16        : out std_logic;
    \-md22\     : out std_logic;
    mf17        : out std_logic;
    \-md21\     : out std_logic;
    mf18        : out std_logic;
    \-md20\     : out std_logic;
    mf19        : out std_logic;
    \-md19\     : out std_logic;
    mf20        : out std_logic;
    \-md18\     : out std_logic;
    mf21        : out std_logic;
    \-md17\     : out std_logic;
    mf22        : out std_logic;
    \-md16\     : out std_logic;
    mf23        : out std_logic;
    \-md7\      : out std_logic;
    mf0         : out std_logic;
    \-md6\      : out std_logic;
    mf1         : out std_logic;
    \-md5\      : out std_logic;
    mf2         : out std_logic;
    \-md4\      : out std_logic;
    mf3         : out std_logic;
    \-md3\      : out std_logic;
    mf4         : out std_logic;
    \-md2\      : out std_logic;
    mf5         : out std_logic;
    \-md1\      : out std_logic;
    mf6         : out std_logic;
    \-md0\      : out std_logic;
    mf7         : out std_logic;
    srcmd       : out std_logic;
    tse2        : in  std_logic;
    \-md15\     : out std_logic;
    mf8         : out std_logic;
    \-md14\     : out std_logic;
    mf9         : out std_logic;
    \-md13\     : out std_logic;
    mf10        : out std_logic;
    \-md12\     : out std_logic;
    mf11        : out std_logic;
    \-md11\     : out std_logic;
    mf12        : out std_logic;
    \-md10\     : out std_logic;
    mf13        : out std_logic;
    \-md9\      : out std_logic;
    mf14        : out std_logic;
    \-md8\      : out std_logic;
    mf15        : out std_logic;
    gnd         : in  std_logic;
    \-mds31\    : in  std_logic;
    \-mds30\    : in  std_logic;
    \-mds29\    : in  std_logic;
    \-mds28\    : in  std_logic;
    mdclk       : out std_logic;
    \-mds27\    : in  std_logic;
    \-mds26\    : in  std_logic;
    \-mds25\    : in  std_logic;
    \-mds24\    : in  std_logic;
    \-mds7\     : in  std_logic;
    \-mds6\     : in  std_logic;
    \-mds5\     : in  std_logic;
    \-mds4\     : in  std_logic;
    \-mds3\     : in  std_logic;
    \-mds2\     : in  std_logic;
    \-mds1\     : in  std_logic;
    \-mds0\     : in  std_logic;
    \-mds23\    : in  std_logic;
    \-mds22\    : in  std_logic;
    \-mds21\    : in  std_logic;
    \-mds20\    : in  std_logic;
    \-mds19\    : in  std_logic;
    \-mds18\    : in  std_logic;
    \-mds17\    : in  std_logic;
    \-mds16\    : in  std_logic;
    destmdr     : out std_logic;
    \-clk2c\    : in  std_logic;
    loadmd      : out std_logic;
    \-loadmd\   : in  std_logic;
    \-destmdr\  : in  std_logic;
    \-mds15\    : in  std_logic;
    \-mds14\    : in  std_logic;
    \-mds13\    : in  std_logic;
    \-mds12\    : in  std_logic;
    \-mds11\    : in  std_logic;
    \-mds10\    : in  std_logic;
    \-mds9\     : in  std_logic;
    \-mds8\     : in  std_logic;
    mdgetspar   : out std_logic;
    \-ignpar\   : in  std_logic;
    mdhaspar    : out std_logic;
    \mempar_in\ : in  std_logic;
    mdpar       : out std_logic;
    \-srcmd\    : in  std_logic);
end;

architecture ttl of cadr4_md is
  signal nc322 : std_logic;
  signal nc323 : std_logic;
  signal nc324 : std_logic;
  signal nc325 : std_logic;
  signal nc326 : std_logic;
  signal nc327 : std_logic;
  signal nc328 : std_logic;
  signal nc329 : std_logic;
  signal nc330 : std_logic;
  signal nc331 : std_logic;
  signal nc332 : std_logic;
  signal nc333 : std_logic;
begin
  md_1a02 : sn74s240 port map(aenb_n => \-mddrive\, ain0 => \-md31\, bout3 => mf24, ain1 => \-md30\, bout2 => mf25, ain2 => \-md29\, bout1 => mf26, ain3 => \-md28\, bout0 => mf27, bin0 => \-md27\, aout3 => mf28, bin1 => \-md26\, aout2 => mf29, bin2 => \-md25\, aout1 => mf30, bin3 => \-md24\, aout0 => mf31, benb_n => \-mddrive\);
  md_1a04 : sn74s240 port map(aenb_n => \-mddrive\, ain0 => \-md23\, bout3 => mf16, ain1 => \-md22\, bout2 => mf17, ain2 => \-md21\, bout1 => mf18, ain3 => \-md20\, bout0 => mf19, bin0 => \-md19\, aout3 => mf20, bin1 => \-md18\, aout2 => mf21, bin2 => \-md17\, aout1 => mf22, bin3 => \-md16\, aout0 => mf23, benb_n => \-mddrive\);
  md_1a05 : sn74s240 port map(aenb_n => \-mddrive\, ain0 => \-md7\, bout3 => mf0, ain1 => \-md6\, bout2 => mf1, ain2 => \-md5\, bout1 => mf2, ain3 => \-md4\, bout0 => mf3, bin0 => \-md3\, aout3 => mf4, bin1 => \-md2\, aout2 => mf5, bin2 => \-md1\, aout1 => mf6, bin3 => \-md0\, aout0 => mf7, benb_n => \-mddrive\);
  md_1a08 : sn74s00 port map(g2b     => srcmd, g2a => tse2, g2q_n => \-mddrive\, g1b => '0', g1a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  md_1a09 : sn74s240 port map(aenb_n => \-mddrive\, ain0 => \-md15\, bout3 => mf8, ain1 => \-md14\, bout2 => mf9, ain2 => \-md13\, bout1 => mf10, ain3 => \-md12\, bout0 => mf11, bin0 => \-md11\, aout3 => mf12, bin1 => \-md10\, aout2 => mf13, bin2 => \-md9\, aout1 => mf14, bin3 => \-md8\, aout0 => mf15, benb_n => \-mddrive\);
  md_1b16 : sn74s374 port map(oenb_n => gnd, o0 => \-md31\, i0 => \-mds31\, i1 => \-mds30\, o1 => \-md30\, o2 => \-md29\, i2 => \-mds29\, i3 => \-mds28\, o3 => \-md28\, clk => mdclk, o4 => \-md27\, i4 => \-mds27\, i5 => \-mds26\, o5 => \-md26\, o6 => \-md25\, i6 => \-mds25\, i7 => \-mds24\, o7 => \-md24\);
  md_1c17 : sn74s374 port map(oenb_n => gnd, o0 => \-md7\, i0 => \-mds7\, i1 => \-mds6\, o1 => \-md6\, o2 => \-md5\, i2 => \-mds5\, i3 => \-mds4\, o3 => \-md4\, clk => mdclk, o4 => \-md3\, i4 => \-mds3\, i5 => \-mds2\, o5 => \-md2\, o6 => \-md1\, i6 => \-mds1\, i7 => \-mds0\, o7 => \-md0\);
  md_1c19 : sn74s374 port map(oenb_n => gnd, o0 => \-md23\, i0 => \-mds23\, i1 => \-mds22\, o1 => \-md22\, o2 => \-md21\, i2 => \-mds21\, i3 => \-mds20\, o3 => \-md20\, clk => mdclk, o4 => \-md19\, i4 => \-mds19\, i5 => \-mds18\, o5 => \-md18\, o6 => \-md17\, i6 => \-mds17\, i7 => \-mds16\, o7 => \-md16\);
  md_1d16 : sn74s51 port map(g2a     => destmdr, g2b => \-clk2c\, g2c => loadmd, g2d => loadmd, g2y => mdclk, g1a => '0', g1c => '0', g1d => '0', g1b => '0');
  md_1d18 : sn74s04 port map(g4q_n   => loadmd, g4a => \-loadmd\, g5q_n => destmdr, g5a => \-destmdr\, g1a => '0', g2a => '0', g3a => '0', g6a => '0');
  md_1d20 : sn74s374 port map(oenb_n => gnd, o0 => \-md15\, i0 => \-mds15\, i1 => \-mds14\, o1 => \-md14\, o2 => \-md13\, i2 => \-mds13\, i3 => \-mds12\, o3 => \-md12\, clk => mdclk, o4 => \-md11\, i4 => \-mds11\, i5 => \-mds10\, o5 => \-md10\, o6 => \-md9\, i6 => \-mds9\, i7 => \-mds8\, o7 => \-md8\);
  md_1e07 : sn74s08 port map(g3q     => mdgetspar, g3a => \-destmdr\, g3b => \-ignpar\, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  md_1e19 : sn74s374 port map(oenb_n => gnd, o0 => nc322, i0 => nc323, i1 => nc324, o1 => nc325, o2 => nc326, i2 => nc327, i3 => nc328, o3 => nc329, clk => mdclk, o4 => nc330, i4 => nc331, i5 => nc332, o5 => nc333, o6 => mdhaspar, i6 => mdgetspar, i7 => \mempar_in\, o7 => mdpar);
  md_2a05 : sn74s04 port map(g2a     => \-srcmd\, g2q_n => srcmd, g1a => '0', g3a => '0', g4a => '0', g5a => '0', g6a => '0');
end architecture;
