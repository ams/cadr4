library ieee;
use ieee.std_logic_1164.all;

-- Dec 14 17:07:30 1980

package icmem_book is
  component cadr_clock1 is
  port (
    \-clock reset b\ : in  std_logic;
    \-hang\          : in  std_logic;
    \-ilong\         : in  std_logic;
    \-tpr0\          : out std_logic;
    \-tpr5\          : out std_logic;
    \-tpr10\         : out std_logic;
    \-tpr15\         : out std_logic;
    \-tpr20\         : out std_logic;
    \-tpr20a\        : out std_logic;
    \-tpr25\         : out std_logic;
    \-tpr40\         : out std_logic;
    \-tpr60\         : out std_logic;
    \-tpr65\         : out std_logic;
    \-tpr70\         : out std_logic;
    \-tpr75\         : out std_logic;
    \-tpr80\         : out std_logic;
    \-tpr80a\        : out std_logic;
    \-tpr85\         : out std_logic;
    \-tpr100\        : out std_logic;
    \-tpr105\        : out std_logic;
    \-tpr110\        : out std_logic;
    \-tpr115\        : out std_logic;
    \-tpr120\        : out std_logic;
    \-tpr120a\       : out std_logic;
    \-tpr125\        : out std_logic;
    \-tpr140\        : out std_logic;
    \-tpr160\        : out std_logic;
    \-tpr180\        : out std_logic;
    \-tpr200\        : out std_logic;
    \-tprend\        : out std_logic;
    \-tpw10\         : out std_logic;
    \-tpw20\         : out std_logic;
    \-tpw25\         : out std_logic;
    \-tpw30\         : out std_logic;
    \-tpw30a\        : out std_logic;
    \-tpw35\         : out std_logic;
    \-tpw40\         : out std_logic;
    \-tpw40a\        : out std_logic;
    \-tpw45\         : out std_logic;
    \-tpw50\         : out std_logic;
    \-tpw55\         : out std_logic;
    \-tpw60\         : out std_logic;
    \-tpw65\         : out std_logic;
    \-tpw70\         : out std_logic;
    \-tpw75\         : out std_logic;
    cyclecompleted   : out std_logic;
    sspeed0          : in  std_logic;
    sspeed1          : in  std_logic;
    tprend           : out std_logic
  );
  end component;
  component cadr_clock2 is
  port (
    \-clk0\          : out std_logic;
    \-clock reset b\ : in  std_logic;
    \-machruna\      : in  std_logic;
    \-mclk0\         : out std_logic;
    \-tpclk\         : out std_logic;
    \-tpr0\          : in  std_logic;
    \-tpr5\          : in  std_logic;
    \-tpr25\         : in  std_logic;
    \-tprend\        : in  std_logic;
    \-tptse\         : out std_logic;
    \-tpw30\         : in  std_logic;
    \-tpw45\         : in  std_logic;
    \-tpw70\         : in  std_logic;
    \-tse1\          : out std_logic;
    \-tse2\          : out std_logic;
    \-tse3\          : out std_logic;
    \-tse4\          : out std_logic;
    \-wp1\           : out std_logic;
    \-wp2\           : out std_logic;
    \-wp3\           : out std_logic;
    \-wp4\           : out std_logic;
    \-wp5\           : out std_logic;
    clk1             : out std_logic;
    clk2             : out std_logic;
    clk3             : out std_logic;
    clk4             : out std_logic;
    clk5             : out std_logic;
    hi1              : in  std_logic;
    machrun          : in  std_logic;
    mclk1            : out std_logic;
    mclk5            : out std_logic;
    mclk7            : out std_logic;
    tpclk            : out std_logic;
    tptse            : out std_logic;
    tpwp             : out std_logic;
    tpwpiram         : out std_logic
  );
  end component;
  component cadr_debug is
  port (
    \-idebug\  : in  std_logic;
    \-lddbirh\ : in  std_logic;
    \-lddbirl\ : in  std_logic;
    \-lddbirm\ : in  std_logic;
    i0         : out std_logic;
    i1         : out std_logic;
    i2         : out std_logic;
    i3         : out std_logic;
    i4         : out std_logic;
    i5         : out std_logic;
    i6         : out std_logic;
    i7         : out std_logic;
    i8         : out std_logic;
    i9         : out std_logic;
    i10        : out std_logic;
    i11        : out std_logic;
    i12        : out std_logic;
    i13        : out std_logic;
    i14        : out std_logic;
    i15        : out std_logic;
    i16        : out std_logic;
    i17        : out std_logic;
    i18        : out std_logic;
    i19        : out std_logic;
    i20        : out std_logic;
    i21        : out std_logic;
    i22        : out std_logic;
    i23        : out std_logic;
    i24        : out std_logic;
    i25        : out std_logic;
    i26        : out std_logic;
    i27        : out std_logic;
    i28        : out std_logic;
    i29        : out std_logic;
    i30        : out std_logic;
    i31        : out std_logic;
    i32        : out std_logic;
    i33        : out std_logic;
    i34        : out std_logic;
    i35        : out std_logic;
    i36        : out std_logic;
    i37        : out std_logic;
    i38        : out std_logic;
    i39        : out std_logic;
    i40        : out std_logic;
    i41        : out std_logic;
    i42        : out std_logic;
    i43        : out std_logic;
    i44        : out std_logic;
    i45        : out std_logic;
    i46        : out std_logic;
    i47        : out std_logic;
    spy0       : in  std_logic;
    spy1       : in  std_logic;
    spy2       : in  std_logic;
    spy3       : in  std_logic;
    spy4       : in  std_logic;
    spy5       : in  std_logic;
    spy6       : in  std_logic;
    spy7       : in  std_logic;
    spy8       : in  std_logic;
    spy9       : in  std_logic;
    spy10      : in  std_logic;
    spy11      : in  std_logic;
    spy12      : in  std_logic;
    spy13      : in  std_logic;
    spy14      : in  std_logic;
    spy15      : in  std_logic
  );
  end component;

--  component cadr_icaps is
--  end component;
  component cadr_ictl is
  port (
    \-ice0a\        : out std_logic;
    \-ice0b\        : out std_logic;
    \-ice0c\        : out std_logic;
    \-ice0d\        : out std_logic;
    \-ice1a\        : out std_logic;
    \-ice1b\        : out std_logic;
    \-ice1c\        : out std_logic;
    \-ice1d\        : out std_logic;
    \-ice2a\        : out std_logic;
    \-ice2b\        : out std_logic;
    \-ice2c\        : out std_logic;
    \-ice2d\        : out std_logic;
    \-ice3a\        : out std_logic;
    \-ice3b\        : out std_logic;
    \-ice3c\        : out std_logic;
    \-ice3d\        : out std_logic;
    \-iwea\         : out std_logic;
    \-iweb\         : out std_logic;
    \-iwec\         : out std_logic;
    \-iwed\         : out std_logic;
    \-iwee\         : out std_logic;
    \-iwef\         : out std_logic;
    \-iweg\         : out std_logic;
    \-iweh\         : out std_logic;
    \-iwei\         : out std_logic;
    \-iwej\         : out std_logic;
    \-iwek\         : out std_logic;
    \-iwel\         : out std_logic;
    \-iwem\         : out std_logic;
    \-iwen\         : out std_logic;
    \-iweo\         : out std_logic;
    \-iwep\         : out std_logic;
    \-iwrited\      : in  std_logic;
    \-iwriteda\     : out std_logic;
    \-pc12b\        : out std_logic;
    \-pc13b\        : out std_logic;
    \-pcb0\         : out std_logic;
    \-pcb1\         : out std_logic;
    \-pcb2\         : out std_logic;
    \-pcb3\         : out std_logic;
    \-pcb4\         : out std_logic;
    \-pcb5\         : out std_logic;
    \-pcb6\         : out std_logic;
    \-pcb7\         : out std_logic;
    \-pcb8\         : out std_logic;
    \-pcb9\         : out std_logic;
    \-pcb10\        : out std_logic;
    \-pcb11\        : out std_logic;
    \-pcc0\         : out std_logic;
    \-pcc1\         : out std_logic;
    \-pcc2\         : out std_logic;
    \-pcc3\         : out std_logic;
    \-pcc4\         : out std_logic;
    \-pcc5\         : out std_logic;
    \-pcc6\         : out std_logic;
    \-pcc7\         : out std_logic;
    \-pcc8\         : out std_logic;
    \-pcc9\         : out std_logic;
    \-pcc10\        : out std_logic;
    \-pcc11\        : out std_logic;
    \-promdisabled\ : out std_logic;
    \-wp5\          : in  std_logic;
    hi1             : in  std_logic;
    idebug          : in  std_logic;
    iwriteda        : out std_logic;
    iwritedb        : out std_logic;
    iwritedc        : out std_logic;
    iwritedd        : out std_logic;
    pc0             : in  std_logic;
    pc1             : in  std_logic;
    pc2             : in  std_logic;
    pc3             : in  std_logic;
    pc4             : in  std_logic;
    pc5             : in  std_logic;
    pc6             : in  std_logic;
    pc7             : in  std_logic;
    pc8             : in  std_logic;
    pc9             : in  std_logic;
    pc10            : in  std_logic;
    pc11            : in  std_logic;
    pc12            : in  std_logic;
    pc13            : in  std_logic;
    promdisabled    : in  std_logic;
    ramdisable      : out std_logic;
    wp5a            : out std_logic;
    wp5b            : out std_logic;
    wp5c            : out std_logic;
    wp5d            : out std_logic
  );
  end component;
  component cadr_iwrpar is
  port (
    iwr0  : in  std_logic;
    iwr1  : in  std_logic;
    iwr2  : in  std_logic;
    iwr3  : in  std_logic;
    iwr4  : in  std_logic;
    iwr5  : in  std_logic;
    iwr6  : in  std_logic;
    iwr7  : in  std_logic;
    iwr8  : in  std_logic;
    iwr9  : in  std_logic;
    iwr10 : in  std_logic;
    iwr11 : in  std_logic;
    iwr12 : in  std_logic;
    iwr13 : in  std_logic;
    iwr14 : in  std_logic;
    iwr15 : in  std_logic;
    iwr16 : in  std_logic;
    iwr17 : in  std_logic;
    iwr18 : in  std_logic;
    iwr19 : in  std_logic;
    iwr20 : in  std_logic;
    iwr21 : in  std_logic;
    iwr22 : in  std_logic;
    iwr23 : in  std_logic;
    iwr24 : in  std_logic;
    iwr25 : in  std_logic;
    iwr26 : in  std_logic;
    iwr27 : in  std_logic;
    iwr28 : in  std_logic;
    iwr29 : in  std_logic;
    iwr30 : in  std_logic;
    iwr31 : in  std_logic;
    iwr32 : in  std_logic;
    iwr33 : in  std_logic;
    iwr34 : in  std_logic;
    iwr35 : in  std_logic;
    iwr36 : in  std_logic;
    iwr37 : in  std_logic;
    iwr38 : in  std_logic;
    iwr39 : in  std_logic;
    iwr40 : in  std_logic;
    iwr41 : in  std_logic;
    iwr42 : in  std_logic;
    iwr43 : in  std_logic;
    iwr44 : in  std_logic;
    iwr45 : in  std_logic;
    iwr46 : in  std_logic;
    iwr47 : in  std_logic;
    iwr48 : out std_logic;
    iwrp1 : out std_logic;
    iwrp2 : out std_logic;
    iwrp3 : out std_logic;
    iwrp4 : out std_logic
  );
  end component;

-- component cadr_mbcpin is
-- end component;

-- component cadr_mcpins is
-- end component;
  component cadr_olord1 is
  port (
    \-boot\          : in  std_logic;
    \-clock reset a\ : in  std_logic;
    \-errhalt\       : in  std_logic;
    \-idebug\        : out std_logic;
    \-ldclk\         : in  std_logic;
    \-ldmode\        : in  std_logic;
    \-ldopc\         : in  std_logic;
    \-ldstat\        : out std_logic;
    \-lpc.hold\      : out std_logic;
    \-machrun\       : out std_logic;
    \-machruna\      : out std_logic;
    \-nop11\         : out std_logic;
    \-opcclk\        : out std_logic;
    \-opcinh\        : out std_logic;
    \-reset\         : in  std_logic;
    \-run\           : out std_logic;
    \-ssdone\        : out std_logic;
    \-stathalt\      : out std_logic;
    \-stc32\         : in  std_logic;
    \-step\          : out std_logic;
    \-tpr60\         : in  std_logic;
    \-wait\          : in  std_logic;
    errstop          : out std_logic;
    idebug           : out std_logic;
    ldstat           : out std_logic;
    \lpc.hold\       : out std_logic;
    machrun          : out std_logic;
    mclk5a           : in  std_logic;
    nop11            : out std_logic;
    opcclk           : out std_logic;
    opcinh           : out std_logic;
    promdisable      : out std_logic;
    promdisabled     : out std_logic;
    run              : out std_logic;
    speed0           : out std_logic;
    speed0a          : out std_logic;
    speed1           : out std_logic;
    speed1a          : out std_logic;
    speedclk         : out std_logic;
    spy0             : in  std_logic;
    spy1             : in  std_logic;
    spy2             : in  std_logic;
    spy3             : in  std_logic;
    spy4             : in  std_logic;
    spy5             : in  std_logic;
    srun             : out std_logic;
    ssdone           : out std_logic;
    sspeed0          : out std_logic;
    sspeed1          : out std_logic;
    sstep            : out std_logic;
    \stat.ovf\       : out std_logic;
    stathenb         : out std_logic;
    statstop         : in  std_logic;
    step             : out std_logic;
    trapenb          : out std_logic
  );
  end component;
  component cadr_olord2 is
  port (
    \-ape\              : out std_logic;
    \-boot1\            : inout std_logic;
    \-boot2\            : out std_logic;
    \-boot\             : out std_logic;
    \-bus.reset\        : out std_logic;
    \-busint.lm.reset\  : in  std_logic;
    \-clk5\             : out std_logic;
    \-clock reset a\    : out std_logic;
    \-clock reset b\    : out std_logic;
    \-dpe\              : out std_logic;
    \-errhalt\          : out std_logic;
    \-halt\             : in  std_logic;
    \-halted\           : out std_logic;
    \-higherr\          : out std_logic;
    \-ipe\              : out std_logic;
    \-ldmode\           : in std_logic;
    \-lowerhighok\      : out std_logic;
    \-mclk5\            : out std_logic;
    \-mempe\            : out std_logic;
    \-mpe\              : out std_logic;
    \-pdlpe\            : out std_logic;
    \-power reset\      : out std_logic;
    \-prog.reset\       : out std_logic;
    \-reset\            : out std_logic;
    \-spe\              : out std_logic;
    \-upperhighok\      : in  std_logic;
    \-v0pe\             : out std_logic;
    \-v1pe\             : out std_logic;
    aparok              : in  std_logic;
    \boot.trap\         : out std_logic;
    \-bus.power.reset\  : out std_logic;
    clk5                : in  std_logic;
    clk5a               : out std_logic;
    dparok              : in  std_logic;
    err                 : out std_logic;
    errstop             : in  std_logic;
    hi1                 : out std_logic;
    hi2                 : out std_logic;
    highok              : out std_logic;
    iparok              : in  std_logic;
    ldmode              : out std_logic;
    mclk5               : in  std_logic;
    mclk5a              : out std_logic;
    memparok            : in  std_logic;
    mmemparok           : in  std_logic;
    pdlparok            : in  std_logic;
    \power reset a\     : out std_logic;
    \prog.boot\         : out std_logic;
    \prog.bus.reset\    : out std_logic;
    reset               : out std_logic;
    spcparok            : in  std_logic;
    spy6                : in  std_logic;
    spy7                : in  std_logic;
    srun                : in  std_logic;
    \stat.ovf\          : in  std_logic;
    statstop            : out std_logic;
    v0parok             : in  std_logic;
    vmoparok            : in  std_logic
  );
  end component;
  component cadr_opcs is
  port (
    \-clk5\   : in  std_logic;
    \-opcinh\ : in  std_logic;
    hi2       : in  std_logic;
    opc0      : out std_logic;
    opc1      : out std_logic;
    opc2      : out std_logic;
    opc3      : out std_logic;
    opc4      : out std_logic;
    opc5      : out std_logic;
    opc6      : out std_logic;
    opc7      : out std_logic;
    opc8      : out std_logic;
    opc9      : out std_logic;
    opc10     : out std_logic;
    opc11     : out std_logic;
    opc12     : out std_logic;
    opc13     : out std_logic;
    opcclk    : in  std_logic;
    opcclka   : out std_logic;
    opcclkb   : out std_logic;
    opcclkc   : out std_logic;
    opcinha   : out std_logic;
    opcinhb   : out std_logic;
    pc0       : in  std_logic;
    pc1       : in  std_logic;
    pc2       : in  std_logic;
    pc3       : in  std_logic;
    pc4       : in  std_logic;
    pc5       : in  std_logic;
    pc6       : in  std_logic;
    pc7       : in  std_logic;
    pc8       : in  std_logic;
    pc9       : in  std_logic;
    pc10      : in  std_logic;
    pc11      : in  std_logic;
    pc12      : in  std_logic;
    pc13      : in  std_logic
  );
  end component;
  component cadr_pctl is
  port (
    \-ape\          : in  std_logic;
    \-dpe\          : in  std_logic;
    \-idebug\       : in  std_logic;
    \-ipe\          : in  std_logic;
    \-iwriteda\     : in  std_logic;
    \-mempe\        : in  std_logic;
    \-mpe\          : in  std_logic;
    \-pdlpe\        : in  std_logic;
    \-promce0\      : out std_logic;
    \-promce1\      : out std_logic;
    \-promdisabled\ : in  std_logic;
    \-promenable\   : out std_logic;
    \-prompc0\      : out std_logic;
    \-prompc1\      : out std_logic;
    \-prompc2\      : out std_logic;
    \-prompc3\      : out std_logic;
    \-prompc4\      : out std_logic;
    \-prompc5\      : out std_logic;
    \-prompc6\      : out std_logic;
    \-prompc7\      : out std_logic;
    \-prompc8\      : out std_logic;
    \-prompc9\      : out std_logic;
    \-spe\          : in  std_logic;
    \-v0pe\         : in  std_logic;
    \-v1pe\         : in  std_logic;
    \bottom.1k\     : out std_logic;
    dpe             : out std_logic;
    hi2             : in  std_logic;
    i46             : out std_logic;
    ipe             : out std_logic;
    pc0             : in  std_logic;
    pc1             : in  std_logic;
    pc2             : in  std_logic;
    pc3             : in  std_logic;
    pc4             : in  std_logic;
    pc5             : in  std_logic;
    pc6             : in  std_logic;
    pc7             : in  std_logic;
    pc8             : in  std_logic;
    pc9             : in  std_logic;
    pc10            : in  std_logic;
    pc11            : in  std_logic;
    pc12            : in  std_logic;
    pc13            : in  std_logic;
    promenable      : out std_logic;
    tilt0           : out std_logic;
    tilt1           : out std_logic
  );
  end component;
  component cadr_prom0 is
  port (
    \-promce0\ : in  std_logic;
    \-prompc0\ : in  std_logic;
    \-prompc1\ : in  std_logic;
    \-prompc2\ : in  std_logic;
    \-prompc3\ : in  std_logic;
    \-prompc4\ : in  std_logic;
    \-prompc5\ : in  std_logic;
    \-prompc6\ : in  std_logic;
    \-prompc7\ : in  std_logic;
    \-prompc8\ : in  std_logic;
    i0         : out std_logic;
    i1         : out std_logic;
    i2         : out std_logic;
    i3         : out std_logic;
    i4         : out std_logic;
    i5         : out std_logic;
    i6         : out std_logic;
    i7         : out std_logic;
    i8         : out std_logic;
    i9         : out std_logic;
    i10        : out std_logic;
    i11        : out std_logic;
    i12        : out std_logic;
    i13        : out std_logic;
    i14        : out std_logic;
    i15        : out std_logic;
    i16        : out std_logic;
    i17        : out std_logic;
    i18        : out std_logic;
    i19        : out std_logic;
    i20        : out std_logic;
    i21        : out std_logic;
    i22        : out std_logic;
    i23        : out std_logic;
    i24        : out std_logic;
    i25        : out std_logic;
    i26        : out std_logic;
    i27        : out std_logic;
    i28        : out std_logic;
    i29        : out std_logic;
    i30        : out std_logic;
    i31        : out std_logic;
    i32        : out std_logic;
    i33        : out std_logic;
    i34        : out std_logic;
    i35        : out std_logic;
    i36        : out std_logic;
    i37        : out std_logic;
    i38        : out std_logic;
    i39        : out std_logic;
    i40        : out std_logic;
    i41        : out std_logic;
    i42        : out std_logic;
    i43        : out std_logic;
    i44        : out std_logic;
    i45        : out std_logic;
    i47        : out std_logic;
    i48        : out std_logic
  );
  end component;
  component cadr_prom1 is
  port (
    \-promce1\ : in  std_logic;
    \-prompc0\ : in  std_logic;
    \-prompc1\ : in  std_logic;
    \-prompc2\ : in  std_logic;
    \-prompc3\ : in  std_logic;
    \-prompc4\ : in  std_logic;
    \-prompc5\ : in  std_logic;
    \-prompc6\ : in  std_logic;
    \-prompc7\ : in  std_logic;
    \-prompc8\ : in  std_logic;
    i0         : out std_logic;
    i1         : out std_logic;
    i2         : out std_logic;
    i3         : out std_logic;
    i4         : out std_logic;
    i5         : out std_logic;
    i6         : out std_logic;
    i7         : out std_logic;
    i8         : out std_logic;
    i9         : out std_logic;
    i10        : out std_logic;
    i11        : out std_logic;
    i12        : out std_logic;
    i13        : out std_logic;
    i14        : out std_logic;
    i15        : out std_logic;
    i16        : out std_logic;
    i17        : out std_logic;
    i18        : out std_logic;
    i19        : out std_logic;
    i20        : out std_logic;
    i21        : out std_logic;
    i22        : out std_logic;
    i23        : out std_logic;
    i24        : out std_logic;
    i25        : out std_logic;
    i26        : out std_logic;
    i27        : out std_logic;
    i28        : out std_logic;
    i29        : out std_logic;
    i30        : out std_logic;
    i31        : out std_logic;
    i32        : out std_logic;
    i33        : out std_logic;
    i34        : out std_logic;
    i35        : out std_logic;
    i36        : out std_logic;
    i37        : out std_logic;
    i38        : out std_logic;
    i39        : out std_logic;
    i40        : out std_logic;
    i41        : out std_logic;
    i42        : out std_logic;
    i43        : out std_logic;
    i44        : out std_logic;
    i45        : out std_logic;
    i47        : out std_logic;
    i48        : out std_logic
  );
  end component;
  component cadr_iram00 is
  port (
    \-ice0a\ : in  std_logic;
    \-iwea\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i0       : out std_logic;
    i1       : out std_logic;
    i2       : out std_logic;
    i3       : out std_logic;
    i4       : out std_logic;
    i5       : out std_logic;
    i6       : out std_logic;
    i7       : out std_logic;
    i8       : out std_logic;
    i9       : out std_logic;
    i10      : out std_logic;
    i11      : out std_logic;
    iwr0     : in  std_logic;
    iwr1     : in  std_logic;
    iwr2     : in  std_logic;
    iwr3     : in  std_logic;
    iwr4     : in  std_logic;
    iwr5     : in  std_logic;
    iwr6     : in  std_logic;
    iwr7     : in  std_logic;
    iwr8     : in  std_logic;
    iwr9     : in  std_logic;
    iwr10    : in  std_logic;
    iwr11    : in  std_logic;
    pc0a     : out std_logic;
    pc1a     : out std_logic;
    pc2a     : out std_logic;
    pc3a     : out std_logic;
    pc4a     : out std_logic;
    pc5a     : out std_logic;
    pc6a     : out std_logic;
    pc7a     : out std_logic;
    pc8a     : out std_logic;
    pc9a     : out std_logic;
    pc10a    : out std_logic;
    pc11a    : out std_logic
  );
  end component;
  component cadr_iram01 is
  port (
    \-ice1a\ : in  std_logic;
    \-iweb\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i0       : out std_logic;
    i1       : out std_logic;
    i2       : out std_logic;
    i3       : out std_logic;
    i4       : out std_logic;
    i5       : out std_logic;
    i6       : out std_logic;
    i7       : out std_logic;
    i8       : out std_logic;
    i9       : out std_logic;
    i10      : out std_logic;
    i11      : out std_logic;
    iwr0     : in  std_logic;
    iwr1     : in  std_logic;
    iwr2     : in  std_logic;
    iwr3     : in  std_logic;
    iwr4     : in  std_logic;
    iwr5     : in  std_logic;
    iwr6     : in  std_logic;
    iwr7     : in  std_logic;
    iwr8     : in  std_logic;
    iwr9     : in  std_logic;
    iwr10    : in  std_logic;
    iwr11    : in  std_logic;
    pc0b     : out std_logic;
    pc1b     : out std_logic;
    pc2b     : out std_logic;
    pc3b     : out std_logic;
    pc4b     : out std_logic;
    pc5b     : out std_logic;
    pc6b     : out std_logic;
    pc7b     : out std_logic;
    pc8b     : out std_logic;
    pc9b     : out std_logic;
    pc10b    : out std_logic;
    pc11b    : out std_logic
  );
  end component;
  component cadr_iram02 is
  port (
    \-ice2a\ : in  std_logic;
    \-iwec\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i0       : out std_logic;
    i1       : out std_logic;
    i2       : out std_logic;
    i3       : out std_logic;
    i4       : out std_logic;
    i5       : out std_logic;
    i6       : out std_logic;
    i7       : out std_logic;
    i8       : out std_logic;
    i9       : out std_logic;
    i10      : out std_logic;
    i11      : out std_logic;
    iwr0     : in  std_logic;
    iwr1     : in  std_logic;
    iwr2     : in  std_logic;
    iwr3     : in  std_logic;
    iwr4     : in  std_logic;
    iwr5     : in  std_logic;
    iwr6     : in  std_logic;
    iwr7     : in  std_logic;
    iwr8     : in  std_logic;
    iwr9     : in  std_logic;
    iwr10    : in  std_logic;
    iwr11    : in  std_logic;
    pc0c     : out std_logic;
    pc1c     : out std_logic;
    pc2c     : out std_logic;
    pc3c     : out std_logic;
    pc4c     : out std_logic;
    pc5c     : out std_logic;
    pc6c     : out std_logic;
    pc7c     : out std_logic;
    pc8c     : out std_logic;
    pc9c     : out std_logic;
    pc10c    : out std_logic;
    pc11c    : out std_logic
  );
  end component;
  component cadr_iram03 is
  port (
    \-ice3a\ : in  std_logic;
    \-iwed\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i0       : out std_logic;
    i1       : out std_logic;
    i2       : out std_logic;
    i3       : out std_logic;
    i4       : out std_logic;
    i5       : out std_logic;
    i6       : out std_logic;
    i7       : out std_logic;
    i8       : out std_logic;
    i9       : out std_logic;
    i10      : out std_logic;
    i11      : out std_logic;
    iwr0     : in  std_logic;
    iwr1     : in  std_logic;
    iwr2     : in  std_logic;
    iwr3     : in  std_logic;
    iwr4     : in  std_logic;
    iwr5     : in  std_logic;
    iwr6     : in  std_logic;
    iwr7     : in  std_logic;
    iwr8     : in  std_logic;
    iwr9     : in  std_logic;
    iwr10    : in  std_logic;
    iwr11    : in  std_logic;
    pc0d     : out std_logic;
    pc1d     : out std_logic;
    pc2d     : out std_logic;
    pc3d     : out std_logic;
    pc4d     : out std_logic;
    pc5d     : out std_logic;
    pc6d     : out std_logic;
    pc7d     : out std_logic;
    pc8d     : out std_logic;
    pc9d     : out std_logic;
    pc10d    : out std_logic;
    pc11d    : out std_logic
  );
  end component;
  component cadr_iram10 is
  port (
    \-ice0b\ : in  std_logic;
    \-iwee\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i12      : out std_logic;
    i13      : out std_logic;
    i14      : out std_logic;
    i15      : out std_logic;
    i16      : out std_logic;
    i17      : out std_logic;
    i18      : out std_logic;
    i19      : out std_logic;
    i20      : out std_logic;
    i21      : out std_logic;
    i22      : out std_logic;
    i23      : out std_logic;
    iwr12    : in  std_logic;
    iwr13    : in  std_logic;
    iwr14    : in  std_logic;
    iwr15    : in  std_logic;
    iwr16    : in  std_logic;
    iwr17    : in  std_logic;
    iwr18    : in  std_logic;
    iwr19    : in  std_logic;
    iwr20    : in  std_logic;
    iwr21    : in  std_logic;
    iwr22    : in  std_logic;
    iwr23    : in  std_logic;
    pc0e     : out std_logic;
    pc1e     : out std_logic;
    pc2e     : out std_logic;
    pc3e     : out std_logic;
    pc4e     : out std_logic;
    pc5e     : out std_logic;
    pc6e     : out std_logic;
    pc7e     : out std_logic;
    pc8e     : out std_logic;
    pc9e     : out std_logic;
    pc10e    : out std_logic;
    pc11e    : out std_logic
  );
  end component;
  component cadr_iram11 is
  port (
    \-ice1b\ : in  std_logic;
    \-iwef\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i12      : out std_logic;
    i13      : out std_logic;
    i14      : out std_logic;
    i15      : out std_logic;
    i16      : out std_logic;
    i17      : out std_logic;
    i18      : out std_logic;
    i19      : out std_logic;
    i20      : out std_logic;
    i21      : out std_logic;
    i22      : out std_logic;
    i23      : out std_logic;
    iwr12    : in  std_logic;
    iwr13    : in  std_logic;
    iwr14    : in  std_logic;
    iwr15    : in  std_logic;
    iwr16    : in  std_logic;
    iwr17    : in  std_logic;
    iwr18    : in  std_logic;
    iwr19    : in  std_logic;
    iwr20    : in  std_logic;
    iwr21    : in  std_logic;
    iwr22    : in  std_logic;
    iwr23    : in  std_logic;
    pc0f     : out std_logic;
    pc1f     : out std_logic;
    pc2f     : out std_logic;
    pc3f     : out std_logic;
    pc4f     : out std_logic;
    pc5f     : out std_logic;
    pc6f     : out std_logic;
    pc7f     : out std_logic;
    pc8f     : out std_logic;
    pc9f     : out std_logic;
    pc10f    : out std_logic;
    pc11f    : out std_logic
  );
  end component;
  component cadr_iram12 is
  port (
    \-ice2b\ : in  std_logic;
    \-iweg\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i12      : out std_logic;
    i13      : out std_logic;
    i14      : out std_logic;
    i15      : out std_logic;
    i16      : out std_logic;
    i17      : out std_logic;
    i18      : out std_logic;
    i19      : out std_logic;
    i20      : out std_logic;
    i21      : out std_logic;
    i22      : out std_logic;
    i23      : out std_logic;
    iwr12    : in  std_logic;
    iwr13    : in  std_logic;
    iwr14    : in  std_logic;
    iwr15    : in  std_logic;
    iwr16    : in  std_logic;
    iwr17    : in  std_logic;
    iwr18    : in  std_logic;
    iwr19    : in  std_logic;
    iwr20    : in  std_logic;
    iwr21    : in  std_logic;
    iwr22    : in  std_logic;
    iwr23    : in  std_logic;
    pc0g     : out std_logic;
    pc1g     : out std_logic;
    pc2g     : out std_logic;
    pc3g     : out std_logic;
    pc4g     : out std_logic;
    pc5g     : out std_logic;
    pc6g     : out std_logic;
    pc7g     : out std_logic;
    pc8g     : out std_logic;
    pc9g     : out std_logic;
    pc10g    : out std_logic;
    pc11g    : out std_logic
  );
  end component;
  component cadr_iram13 is
  port (
    \-ice3b\ : in  std_logic;
    \-iweh\  : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    i12      : out std_logic;
    i13      : out std_logic;
    i14      : out std_logic;
    i15      : out std_logic;
    i16      : out std_logic;
    i17      : out std_logic;
    i18      : out std_logic;
    i19      : out std_logic;
    i20      : out std_logic;
    i21      : out std_logic;
    i22      : out std_logic;
    i23      : out std_logic;
    iwr12    : in  std_logic;
    iwr13    : in  std_logic;
    iwr14    : in  std_logic;
    iwr15    : in  std_logic;
    iwr16    : in  std_logic;
    iwr17    : in  std_logic;
    iwr18    : in  std_logic;
    iwr19    : in  std_logic;
    iwr20    : in  std_logic;
    iwr21    : in  std_logic;
    iwr22    : in  std_logic;
    iwr23    : in  std_logic;
    pc0h     : out std_logic;
    pc1h     : out std_logic;
    pc2h     : out std_logic;
    pc3h     : out std_logic;
    pc4h     : out std_logic;
    pc5h     : out std_logic;
    pc6h     : out std_logic;
    pc7h     : out std_logic;
    pc8h     : out std_logic;
    pc9h     : out std_logic;
    pc10h    : out std_logic;
    pc11h    : out std_logic
  );
  end component;
  component cadr_iram20 is
  port (
    \-ice0c\ : in  std_logic;
    \-iwei\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i24      : out std_logic;
    i25      : out std_logic;
    i26      : out std_logic;
    i27      : out std_logic;
    i28      : out std_logic;
    i29      : out std_logic;
    i30      : out std_logic;
    i31      : out std_logic;
    i32      : out std_logic;
    i33      : out std_logic;
    i34      : out std_logic;
    i35      : out std_logic;
    iwr24    : in  std_logic;
    iwr25    : in  std_logic;
    iwr26    : in  std_logic;
    iwr27    : in  std_logic;
    iwr28    : in  std_logic;
    iwr29    : in  std_logic;
    iwr30    : in  std_logic;
    iwr31    : in  std_logic;
    iwr32    : in  std_logic;
    iwr33    : in  std_logic;
    iwr34    : in  std_logic;
    iwr35    : in  std_logic;
    pc0i     : out std_logic;
    pc1i     : out std_logic;
    pc2i     : out std_logic;
    pc3i     : out std_logic;
    pc4i     : out std_logic;
    pc5i     : out std_logic;
    pc6i     : out std_logic;
    pc7i     : out std_logic;
    pc8i     : out std_logic;
    pc9i     : out std_logic;
    pc10i    : out std_logic;
    pc11i    : out std_logic
  );
  end component;
  component cadr_iram21 is
  port (
    \-ice1c\ : in  std_logic;
    \-iwej\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i24      : out std_logic;
    i25      : out std_logic;
    i26      : out std_logic;
    i27      : out std_logic;
    i28      : out std_logic;
    i29      : out std_logic;
    i30      : out std_logic;
    i31      : out std_logic;
    i32      : out std_logic;
    i33      : out std_logic;
    i34      : out std_logic;
    i35      : out std_logic;
    iwr24    : in  std_logic;
    iwr25    : in  std_logic;
    iwr26    : in  std_logic;
    iwr27    : in  std_logic;
    iwr28    : in  std_logic;
    iwr29    : in  std_logic;
    iwr30    : in  std_logic;
    iwr31    : in  std_logic;
    iwr32    : in  std_logic;
    iwr33    : in  std_logic;
    iwr34    : in  std_logic;
    iwr35    : in  std_logic;
    pc0j     : out std_logic;
    pc1j     : out std_logic;
    pc2j     : out std_logic;
    pc3j     : out std_logic;
    pc4j     : out std_logic;
    pc5j     : out std_logic;
    pc6j     : out std_logic;
    pc7j     : out std_logic;
    pc8j     : out std_logic;
    pc9j     : out std_logic;
    pc10j    : out std_logic;
    pc11j    : out std_logic
  );
  end component;
  component cadr_iram22 is
  port (
    \-ice2c\ : in  std_logic;
    \-iwek\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i24      : out std_logic;
    i25      : out std_logic;
    i26      : out std_logic;
    i27      : out std_logic;
    i28      : out std_logic;
    i29      : out std_logic;
    i30      : out std_logic;
    i31      : out std_logic;
    i32      : out std_logic;
    i33      : out std_logic;
    i34      : out std_logic;
    i35      : out std_logic;
    iwr24    : in  std_logic;
    iwr25    : in  std_logic;
    iwr26    : in  std_logic;
    iwr27    : in  std_logic;
    iwr28    : in  std_logic;
    iwr29    : in  std_logic;
    iwr30    : in  std_logic;
    iwr31    : in  std_logic;
    iwr32    : in  std_logic;
    iwr33    : in  std_logic;
    iwr34    : in  std_logic;
    iwr35    : in  std_logic;
    pc0k     : out std_logic;
    pc1k     : out std_logic;
    pc2k     : out std_logic;
    pc3k     : out std_logic;
    pc4k     : out std_logic;
    pc5k     : out std_logic;
    pc6k     : out std_logic;
    pc7k     : out std_logic;
    pc8k     : out std_logic;
    pc9k     : out std_logic;
    pc10k    : out std_logic;
    pc11k    : out std_logic
  );
  end component;
  component cadr_iram23 is
  port (
    \-ice3c\ : in  std_logic;
    \-iwel\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i24      : out std_logic;
    i25      : out std_logic;
    i26      : out std_logic;
    i27      : out std_logic;
    i28      : out std_logic;
    i29      : out std_logic;
    i30      : out std_logic;
    i31      : out std_logic;
    i32      : out std_logic;
    i33      : out std_logic;
    i34      : out std_logic;
    i35      : out std_logic;
    iwr24    : in  std_logic;
    iwr25    : in  std_logic;
    iwr26    : in  std_logic;
    iwr27    : in  std_logic;
    iwr28    : in  std_logic;
    iwr29    : in  std_logic;
    iwr30    : in  std_logic;
    iwr31    : in  std_logic;
    iwr32    : in  std_logic;
    iwr33    : in  std_logic;
    iwr34    : in  std_logic;
    iwr35    : in  std_logic;
    pc0l     : out std_logic;
    pc1l     : out std_logic;
    pc2l     : out std_logic;
    pc3l     : out std_logic;
    pc4l     : out std_logic;
    pc5l     : out std_logic;
    pc6l     : out std_logic;
    pc7l     : out std_logic;
    pc8l     : out std_logic;
    pc9l     : out std_logic;
    pc10l    : out std_logic;
    pc11l    : out std_logic
  );
  end component;
  component cadr_iram30 is
  port (
    \-ice0d\ : in  std_logic;
    \-iwem\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i36      : out std_logic;
    i37      : out std_logic;
    i38      : out std_logic;
    i39      : out std_logic;
    i40      : out std_logic;
    i41      : out std_logic;
    i42      : out std_logic;
    i43      : out std_logic;
    i44      : out std_logic;
    i45      : out std_logic;
    i46      : out std_logic;
    i47      : out std_logic;
    i48      : out std_logic;
    iwr36    : in  std_logic;
    iwr37    : in  std_logic;
    iwr38    : in  std_logic;
    iwr39    : in  std_logic;
    iwr40    : in  std_logic;
    iwr41    : in  std_logic;
    iwr42    : in  std_logic;
    iwr43    : in  std_logic;
    iwr44    : in  std_logic;
    iwr45    : in  std_logic;
    iwr46    : in  std_logic;
    iwr47    : in  std_logic;
    iwr48    : in  std_logic;
    pc0m     : out std_logic;
    pc1m     : out std_logic;
    pc2m     : out std_logic;
    pc3m     : out std_logic;
    pc4m     : out std_logic;
    pc5m     : out std_logic;
    pc6m     : out std_logic;
    pc7m     : out std_logic;
    pc8m     : out std_logic;
    pc9m     : out std_logic;
    pc10m    : out std_logic;
    pc11m    : out std_logic
  );
  end component;
  component cadr_iram31 is
  port (
    \-ice1d\ : in  std_logic;
    \-iwen\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i36      : out std_logic;
    i37      : out std_logic;
    i38      : out std_logic;
    i39      : out std_logic;
    i40      : out std_logic;
    i41      : out std_logic;
    i42      : out std_logic;
    i43      : out std_logic;
    i44      : out std_logic;
    i45      : out std_logic;
    i46      : out std_logic;
    i47      : out std_logic;
    i48      : out std_logic;
    iwr36    : in  std_logic;
    iwr37    : in  std_logic;
    iwr38    : in  std_logic;
    iwr39    : in  std_logic;
    iwr40    : in  std_logic;
    iwr41    : in  std_logic;
    iwr42    : in  std_logic;
    iwr43    : in  std_logic;
    iwr44    : in  std_logic;
    iwr45    : in  std_logic;
    iwr46    : in  std_logic;
    iwr47    : in  std_logic;
    iwr48    : in  std_logic;
    pc0n     : out std_logic;
    pc1n     : out std_logic;
    pc2n     : out std_logic;
    pc3n     : out std_logic;
    pc4n     : out std_logic;
    pc5n     : out std_logic;
    pc6n     : out std_logic;
    pc7n     : out std_logic;
    pc8n     : out std_logic;
    pc9n     : out std_logic;
    pc10n    : out std_logic;
    pc11n    : out std_logic
  );
  end component;
  component cadr_iram32 is
  port (
    \-ice2d\ : in  std_logic;
    \-iweo\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i36      : out std_logic;
    i37      : out std_logic;
    i38      : out std_logic;
    i39      : out std_logic;
    i40      : out std_logic;
    i41      : out std_logic;
    i42      : out std_logic;
    i43      : out std_logic;
    i44      : out std_logic;
    i45      : out std_logic;
    i46      : out std_logic;
    i47      : out std_logic;
    i48      : out std_logic;
    iwr36    : in  std_logic;
    iwr37    : in  std_logic;
    iwr38    : in  std_logic;
    iwr39    : in  std_logic;
    iwr40    : in  std_logic;
    iwr41    : in  std_logic;
    iwr42    : in  std_logic;
    iwr43    : in  std_logic;
    iwr44    : in  std_logic;
    iwr45    : in  std_logic;
    iwr46    : in  std_logic;
    iwr47    : in  std_logic;
    iwr48    : in  std_logic;
    pc0o     : out std_logic;
    pc1o     : out std_logic;
    pc2o     : out std_logic;
    pc3o     : out std_logic;
    pc4o     : out std_logic;
    pc5o     : out std_logic;
    pc6o     : out std_logic;
    pc7o     : out std_logic;
    pc8o     : out std_logic;
    pc9o     : out std_logic;
    pc10o    : out std_logic;
    pc11o    : out std_logic
  );
  end component;
  component cadr_iram33 is
  port (
    \-ice3d\ : in  std_logic;
    \-iwep\  : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    i36      : out std_logic;
    i37      : out std_logic;
    i38      : out std_logic;
    i39      : out std_logic;
    i40      : out std_logic;
    i41      : out std_logic;
    i42      : out std_logic;
    i43      : out std_logic;
    i44      : out std_logic;
    i45      : out std_logic;
    i46      : out std_logic;
    i47      : out std_logic;
    i48      : out std_logic;
    iwr36    : in  std_logic;
    iwr37    : in  std_logic;
    iwr38    : in  std_logic;
    iwr39    : in  std_logic;
    iwr40    : in  std_logic;
    iwr41    : in  std_logic;
    iwr42    : in  std_logic;
    iwr43    : in  std_logic;
    iwr44    : in  std_logic;
    iwr45    : in  std_logic;
    iwr46    : in  std_logic;
    iwr47    : in  std_logic;
    iwr48    : in  std_logic;
    pc0p     : out std_logic;
    pc1p     : out std_logic;
    pc2p     : out std_logic;
    pc3p     : out std_logic;
    pc4p     : out std_logic;
    pc5p     : out std_logic;
    pc6p     : out std_logic;
    pc7p     : out std_logic;
    pc8p     : out std_logic;
    pc9p     : out std_logic;
    pc10p    : out std_logic;
    pc11p    : out std_logic
  );
  end component;
  component cadr_spy0 is
  port (
    \-dbread\    : in  std_logic;
    \-dbwrite\   : in  std_logic;
    \-ldclk\     : out std_logic;
    \-lddbirh\   : out std_logic;
    \-lddbirl\   : out std_logic;
    \-lddbirm\   : out std_logic;
    \-ldmode\    : out std_logic;
    \-ldopc\     : out std_logic;
    \-spy.ah\    : out std_logic;
    \-spy.al\    : out std_logic;
    \-spy.flag1\ : out std_logic;
    \-spy.flag2\ : out std_logic;
    \-spy.irh\   : out std_logic;
    \-spy.irl\   : out std_logic;
    \-spy.irm\   : out std_logic;
    \-spy.mh\    : out std_logic;
    \-spy.ml\    : out std_logic;
    \-spy.obh\   : out std_logic;
    \-spy.obl\   : out std_logic;
    \-spy.opc\   : out std_logic;
    \-spy.pc\    : out std_logic;
    \-spy.sth\   : out std_logic;
    \-spy.stl\   : out std_logic;
    eadr0        : in  std_logic;
    eadr1        : in  std_logic;
    eadr2        : in  std_logic;
    eadr3        : in  std_logic;
    hi1          : in  std_logic
  );
  end component;
  component cadr_spy4 is
  port (
    \-ape\       : in  std_logic;
    \-dpe\       : in  std_logic;
    \-higherr\   : in  std_logic;
    \-ipe\       : in  std_logic;
    \-mempe\     : in  std_logic;
    \-mpe\       : in  std_logic;
    \-pdlpe\     : in  std_logic;
    \-spe\       : in  std_logic;
    \-spy.flag1\ : out std_logic;
    \-spy.opc\   : in  std_logic;
    \-spy.pc\    : in  std_logic;
    \-stathalt\  : in  std_logic;
    \-v0pe\      : in  std_logic;
    \-v1pe\      : in  std_logic;
    \-wait\      : in  std_logic;
    err          : in  std_logic;
    opc0         : in  std_logic;
    opc1         : in  std_logic;
    opc2         : in  std_logic;
    opc3         : in  std_logic;
    opc4         : in  std_logic;
    opc5         : in  std_logic;
    opc6         : in  std_logic;
    opc7         : in  std_logic;
    opc8         : in  std_logic;
    opc9         : in  std_logic;
    opc10        : in  std_logic;
    opc11        : in  std_logic;
    opc12        : in  std_logic;
    opc13        : in  std_logic;
    pc0          : in  std_logic;
    pc1          : in  std_logic;
    pc2          : in  std_logic;
    pc3          : in  std_logic;
    pc4          : in  std_logic;
    pc5          : in  std_logic;
    pc6          : in  std_logic;
    pc7          : in  std_logic;
    pc8          : in  std_logic;
    pc9          : in  std_logic;
    pc10         : in  std_logic;
    pc11         : in  std_logic;
    pc12         : in  std_logic;
    pc13         : in  std_logic;
    promdisable  : in  std_logic;
    spy0         : out std_logic;
    spy1         : out std_logic;
    spy2         : out std_logic;
    spy3         : out std_logic;
    spy4         : out std_logic;
    spy5         : out std_logic;
    spy6         : out std_logic;
    spy7         : out std_logic;
    spy8         : out std_logic;
    spy9         : out std_logic;
    spy10        : out std_logic;
    spy11        : out std_logic;
    spy12        : out std_logic;
    spy13        : out std_logic;
    spy14        : out std_logic;
    spy15        : out std_logic;
    srun         : in  std_logic;
    ssdone       : in  std_logic
  );
  end component;
  component cadr_stat is
  port (
    \-ldstat\  : in  std_logic;
    \-spy.sth\ : in  std_logic;
    \-spy.stl\ : in  std_logic;
    \-statbit\ : in  std_logic;
    \-stc4\    : out std_logic;
    \-stc8\    : out std_logic;
    \-stc12\   : out std_logic;
    \-stc16\   : out std_logic;
    \-stc20\   : out std_logic;
    \-stc24\   : out std_logic;
    \-stc28\   : out std_logic;
    \-stc32\   : out std_logic;
    clk5a      : in  std_logic;
    hi1        : in  std_logic;
    iwr0       : in  std_logic;
    iwr1       : in  std_logic;
    iwr2       : in  std_logic;
    iwr3       : in  std_logic;
    iwr4       : in  std_logic;
    iwr5       : in  std_logic;
    iwr6       : in  std_logic;
    iwr7       : in  std_logic;
    iwr8       : in  std_logic;
    iwr9       : in  std_logic;
    iwr10      : in  std_logic;
    iwr11      : in  std_logic;
    iwr12      : in  std_logic;
    iwr13      : in  std_logic;
    iwr14      : in  std_logic;
    iwr15      : in  std_logic;
    iwr16      : in  std_logic;
    iwr17      : in  std_logic;
    iwr18      : in  std_logic;
    iwr19      : in  std_logic;
    iwr20      : in  std_logic;
    iwr21      : in  std_logic;
    iwr22      : in  std_logic;
    iwr23      : in  std_logic;
    iwr24      : in  std_logic;
    iwr25      : in  std_logic;
    iwr26      : in  std_logic;
    iwr27      : in  std_logic;
    iwr28      : in  std_logic;
    iwr29      : in  std_logic;
    iwr30      : in  std_logic;
    iwr31      : in  std_logic;
    spy0       : out std_logic;
    spy1       : out std_logic;
    spy2       : out std_logic;
    spy3       : out std_logic;
    spy4       : out std_logic;
    spy5       : out std_logic;
    spy6       : out std_logic;
    spy7       : out std_logic;
    spy8       : out std_logic;
    spy9       : out std_logic;
    spy10      : out std_logic;
    spy11      : out std_logic;
    spy12      : out std_logic;
    spy13      : out std_logic;
    spy14      : out std_logic;
    spy15      : out std_logic;
    st0        : out std_logic;
    st1        : out std_logic;
    st2        : out std_logic;
    st3        : out std_logic;
    st4        : out std_logic;
    st5        : out std_logic;
    st6        : out std_logic;
    st7        : out std_logic;
    st8        : out std_logic;
    st9        : out std_logic;
    st10       : out std_logic;
    st11       : out std_logic;
    st12       : out std_logic;
    st13       : out std_logic;
    st14       : out std_logic;
    st15       : out std_logic;
    st16       : out std_logic;
    st17       : out std_logic;
    st18       : out std_logic;
    st19       : out std_logic;
    st20       : out std_logic;
    st21       : out std_logic;
    st22       : out std_logic;
    st23       : out std_logic;
    st24       : out std_logic;
    st25       : out std_logic;
    st26       : out std_logic;
    st27       : out std_logic;
    st28       : out std_logic;
    st29       : out std_logic;
    st30       : out std_logic;
    st31       : out std_logic
  );
  end component;

end package;
