library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn7428_tb is
end sn7428_tb;

architecture testbench of sn7428_tb is

begin

--  uut : sn7428 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
