-- CADR1_XAPAR
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_xapar is
  port (
    \xao 0\ : in std_logic;
    \xao 1\ : in std_logic;
    \xao 10\ : in std_logic;
    \xao 11\ : in std_logic;
    \xao 12\ : in std_logic;
    \xao 13\ : in std_logic;
    \xao 14\ : in std_logic;
    \xao 15\ : in std_logic;
    \xao 16\ : in std_logic;
    \xao 17\ : in std_logic;
    \xao 18\ : in std_logic;
    \xao 19\ : in std_logic;
    \xao 2\ : in std_logic;
    \xao 20\ : in std_logic;
    \xao 21\ : in std_logic;
    \xao 3\ : in std_logic;
    \xao 4\ : in std_logic;
    \xao 5\ : in std_logic;
    \xao 6\ : in std_logic;
    \xao 7\ : in std_logic;
    \xao 8\ : in std_logic;
    \xao 9\ : in std_logic;
    \xao par even\ : out std_logic;
    \xao par odd\ : out std_logic
  );
end entity;
