library ieee;
use ieee.std_logic_1164.all;

package set is
  component alu_set is
      -- internal signals: aluf0a aluf0b aluf1a aluf1b aluf2a 
      -- internal signals: aluf2b aluf3a aluf3b alumode \-cin0\ 
      -- internal signals: \-cin4\ \-cin8\ \-cin12\ \-cin16\ \-cin20\ 
      -- internal signals: \-cin24\ \-cin28\ \-cin32\ xout3 xout7 
      -- internal signals: xout11 xout19 xout23 xout27 yout3 
      -- internal signals: yout7 yout11 yout19 yout23 yout27 
    port (
      a0: in std_logic;
      a1: in std_logic;
      a2: in std_logic;
      a3: in std_logic;
      a4: in std_logic;
      a5: in std_logic;
      a6: in std_logic;
      a7: in std_logic;
      a8: in std_logic;
      a9: in std_logic;
      a10: in std_logic;
      a11: in std_logic;
      a13: in std_logic;
      a14: in std_logic;
      a15: in std_logic;
      a16: in std_logic;
      a17: in std_logic;
      a18: in std_logic;
      a19: in std_logic;
      a20: in std_logic;
      a21: in std_logic;
      a22: in std_logic;
      a23: in std_logic;
      a24: in std_logic;
      a25: in std_logic;
      a26: in std_logic;
      a27: in std_logic;
      a28: in std_logic;
      a29: in std_logic;
      a30: in std_logic;
      a31a: in std_logic;
      a31b: in std_logic;
      \-div\: in std_logic;
      hi12: in std_logic;
      ir0: in std_logic;
      ir1: in std_logic;
      ir2: in std_logic;
      ir3: in std_logic;
      ir4: in std_logic;
      ir5: in std_logic;
      ir6: in std_logic;
      ir7: in std_logic;
      \-ir12\: in std_logic;
      \-ir13\: in std_logic;
      \-iralu\: in std_logic;
      irjump: in std_logic;
      \-irjump\: in std_logic;
      m0: in std_logic;
      m1: in std_logic;
      m2: in std_logic;
      m3: in std_logic;
      m4: in std_logic;
      m5: in std_logic;
      m6: in std_logic;
      m7: in std_logic;
      m8: in std_logic;
      m9: in std_logic;
      m10: in std_logic;
      m11: in std_logic;
      m12: in std_logic;
      m13: in std_logic;
      m14: in std_logic;
      m15: in std_logic;
      m16: in std_logic;
      m17: in std_logic;
      m18: in std_logic;
      m19: in std_logic;
      m20: in std_logic;
      m21: in std_logic;
      m22: in std_logic;
      m23: in std_logic;
      m24: in std_logic;
      m25: in std_logic;
      m26: in std_logic;
      m27: in std_logic;
      m28: in std_logic;
      m29: in std_logic;
      m30: in std_logic;
      m31: in std_logic;
      \-mul\: in std_logic;
      q0: in std_logic;
      a12: out std_logic;
      \a=m\: out std_logic;
      alu0: out std_logic;
      alu1: out std_logic;
      alu2: out std_logic;
      alu3: out std_logic;
      alu4: out std_logic;
      alu5: out std_logic;
      alu6: out std_logic;
      alu7: out std_logic;
      alu8: out std_logic;
      alu9: out std_logic;
      alu10: out std_logic;
      alu11: out std_logic;
      alu12: out std_logic;
      alu13: out std_logic;
      alu14: out std_logic;
      alu15: out std_logic;
      alu16: out std_logic;
      alu17: out std_logic;
      alu18: out std_logic;
      alu19: out std_logic;
      alu20: out std_logic;
      alu21: out std_logic;
      alu22: out std_logic;
      alu23: out std_logic;
      alu24: out std_logic;
      alu25: out std_logic;
      alu26: out std_logic;
      alu27: out std_logic;
      alu28: out std_logic;
      alu29: out std_logic;
      alu30: out std_logic;
      alu31: out std_logic;
      alu32: out std_logic;
      \-ir0\: out std_logic;
      \-ir1\: out std_logic;
      \-ir2\: out std_logic;
      \-ir3\: out std_logic;
      \-ir4\: out std_logic;
      osel0a: out std_logic;
      osel0b: out std_logic;
      osel1a: out std_logic;
      osel1b: out std_logic
    );
  end component;
  component amem_set is
      -- internal signals: \-aadr0a\ \-aadr0b\ \-aadr1a\ \-aadr1b\ \-aadr2a\ 
      -- internal signals: \-aadr2b\ \-aadr3a\ \-aadr3b\ \-aadr4a\ \-aadr4b\ 
      -- internal signals: \-aadr5a\ \-aadr5b\ \-aadr6a\ \-aadr6b\ \-aadr7a\ 
      -- internal signals: \-aadr7b\ \-aadr8a\ \-aadr8b\ \-aadr9a\ \-aadr9b\ 
      -- internal signals: amem0 amem1 amem2 amem3 amem4 
      -- internal signals: amem5 amem6 amem7 amem8 amem9 
      -- internal signals: amem10 amem11 amem12 amem13 amem14 
      -- internal signals: amem15 amem16 amem17 amem18 amem19 
      -- internal signals: amem20 amem21 amem22 amem23 amem24 
      -- internal signals: amem25 amem26 amem27 amem28 amem29 
      -- internal signals: amem30 amem31 \-amemenb\ amemparity apassenb 
      -- internal signals: \-apassenb\ \-awpa\ \-awpb\ \-awpc\ 
    port (
      clk3d: in std_logic;
      clk3e: in std_logic;
      dest: in std_logic;
      destm: in std_logic;
      hi3: in std_logic;
      hi5: in std_logic;
      ir14: in std_logic;
      ir15: in std_logic;
      ir16: in std_logic;
      ir17: in std_logic;
      ir18: in std_logic;
      ir19: in std_logic;
      ir20: in std_logic;
      ir21: in std_logic;
      ir22: in std_logic;
      ir23: in std_logic;
      ir32: in std_logic;
      ir33: in std_logic;
      ir34: in std_logic;
      ir35: in std_logic;
      ir36: in std_logic;
      ir37: in std_logic;
      ir38: in std_logic;
      ir39: in std_logic;
      ir40: in std_logic;
      ir41: in std_logic;
      l0: in std_logic;
      l1: in std_logic;
      l2: in std_logic;
      l3: in std_logic;
      l4: in std_logic;
      l5: in std_logic;
      l6: in std_logic;
      l7: in std_logic;
      l8: in std_logic;
      l9: in std_logic;
      l10: in std_logic;
      l11: in std_logic;
      l12: in std_logic;
      l13: in std_logic;
      l14: in std_logic;
      l15: in std_logic;
      l16: in std_logic;
      l17: in std_logic;
      l18: in std_logic;
      l19: in std_logic;
      l20: in std_logic;
      l21: in std_logic;
      l22: in std_logic;
      l23: in std_logic;
      l24: in std_logic;
      l25: in std_logic;
      l26: in std_logic;
      l27: in std_logic;
      l28: in std_logic;
      l29: in std_logic;
      l30: in std_logic;
      l31: in std_logic;
      lparity: in std_logic;
      \-reset\: in std_logic;
      tse3a: in std_logic;
      tse4a: in std_logic;
      wp3a: in std_logic;
      a0: out std_logic;
      a1: out std_logic;
      a2: out std_logic;
      a3: out std_logic;
      a4: out std_logic;
      a5: out std_logic;
      a6: out std_logic;
      a7: out std_logic;
      a8: out std_logic;
      a9: out std_logic;
      a10: out std_logic;
      a11: out std_logic;
      a12: out std_logic;
      a13: out std_logic;
      a14: out std_logic;
      a15: out std_logic;
      a16: out std_logic;
      a17: out std_logic;
      a18: out std_logic;
      a19: out std_logic;
      a20: out std_logic;
      a21: out std_logic;
      a22: out std_logic;
      a23: out std_logic;
      a24: out std_logic;
      a25: out std_logic;
      a26: out std_logic;
      a27: out std_logic;
      a28: out std_logic;
      a29: out std_logic;
      a30: out std_logic;
      a31a: out std_logic;
      a31b: out std_logic;
      aparity: out std_logic;
      destmd: out std_logic;
      wadr0: out std_logic;
      wadr1: out std_logic;
      wadr2: out std_logic;
      wadr3: out std_logic;
      wadr4: out std_logic
    );
  end component;
  component ampar_set is

    port (
      a0: in std_logic;
      a1: in std_logic;
      a2: in std_logic;
      a3: in std_logic;
      a4: in std_logic;
      a5: in std_logic;
      a6: in std_logic;
      a7: in std_logic;
      a8: in std_logic;
      a9: in std_logic;
      a10: in std_logic;
      a11: in std_logic;
      a12: in std_logic;
      a13: in std_logic;
      a14: in std_logic;
      a15: in std_logic;
      a16: in std_logic;
      a17: in std_logic;
      a18: in std_logic;
      a19: in std_logic;
      a20: in std_logic;
      a21: in std_logic;
      a22: in std_logic;
      a23: in std_logic;
      a24: in std_logic;
      a25: in std_logic;
      a26: in std_logic;
      a27: in std_logic;
      a28: in std_logic;
      a29: in std_logic;
      a30: in std_logic;
      a31b: in std_logic;
      aparity: in std_logic;
      m0: in std_logic;
      m1: in std_logic;
      m2: in std_logic;
      m3: in std_logic;
      m4: in std_logic;
      m5: in std_logic;
      m6: in std_logic;
      m7: in std_logic;
      m8: in std_logic;
      m9: in std_logic;
      m10: in std_logic;
      m11: in std_logic;
      m12: in std_logic;
      m13: in std_logic;
      m14: in std_logic;
      m15: in std_logic;
      m16: in std_logic;
      m17: in std_logic;
      m18: in std_logic;
      m19: in std_logic;
      m20: in std_logic;
      m21: in std_logic;
      m22: in std_logic;
      m23: in std_logic;
      m24: in std_logic;
      m25: in std_logic;
      m26: in std_logic;
      m27: in std_logic;
      m28: in std_logic;
      m29: in std_logic;
      m30: in std_logic;
      m31: in std_logic;
      mparity: in std_logic;
      pdlenb: in std_logic;
      srcm: in std_logic;
      aparok: out std_logic;
      mmemparok: out std_logic;
      pdlparok: out std_logic
    );
  end component;
  component clock_set is
      -- internal signals: clk1 clk2 clk3 clk4 mclk1 
      -- internal signals: \-tpr0\ \-tpr5\ \-tpr25\ \-tprend\ \-tpw30\ 
      -- internal signals: \-tpw45\ \-tpw70\ \-tse1\ \-tse2\ \-tse3\ 
      -- internal signals: \-tse4\ \-wp1\ \-wp2\ \-wp3\ \-wp4\ 
    port (
      \-clock reset b\: in std_logic;
      \-hang\: in std_logic;
      hi1: in std_logic;
      hi2: in std_logic;
      hi3: in std_logic;
      hi4: in std_logic;
      hi5: in std_logic;
      hi6: in std_logic;
      hi7: in std_logic;
      hi8: in std_logic;
      hi9: in std_logic;
      hi10: in std_logic;
      hi11: in std_logic;
      hi12: in std_logic;
      \-ilong\: in std_logic;
      lcry3: in std_logic;
      machrun: in std_logic;
      \-machruna\: in std_logic;
      reset: in std_logic;
      \-srcpdlidx\: in std_logic;
      \-srcpdlptr\: in std_logic;
      sspeed0: in std_logic;
      sspeed1: in std_logic;
      clk5: out std_logic;
      clk1a: out std_logic;
      clk2a: out std_logic;
      clk2b: out std_logic;
      clk2c: out std_logic;
      clk3a: out std_logic;
      clk3b: out std_logic;
      clk3c: out std_logic;
      clk3d: out std_logic;
      clk3e: out std_logic;
      clk3f: out std_logic;
      clk4a: out std_logic;
      clk4b: out std_logic;
      clk4c: out std_logic;
      clk4d: out std_logic;
      clk4e: out std_logic;
      clk4f: out std_logic;
      \-clk2c\: out std_logic;
      \-clk3g\: out std_logic;
      \-clk4e\: out std_logic;
      \-lcry3\: out std_logic;
      mclk5: out std_logic;
      mclk1a: out std_logic;
      \-reset\: out std_logic;
      srcpdlidx: out std_logic;
      srcpdlptr: out std_logic;
      \-tpr60\: out std_logic;
      tse2: out std_logic;
      tse1a: out std_logic;
      tse1b: out std_logic;
      tse3a: out std_logic;
      tse4a: out std_logic;
      tse4b: out std_logic;
      \-upperhighok\: out std_logic;
      wp2: out std_logic;
      wp1a: out std_logic;
      wp1b: out std_logic;
      wp3a: out std_logic;
      wp4a: out std_logic;
      wp4b: out std_logic;
      wp4c: out std_logic;
      \-wp5\: out std_logic
    );
  end component;
  component decode_set is

    port (
      hi5: in std_logic;
      \-idebug\: in std_logic;
      ir3: in std_logic;
      ir4: in std_logic;
      ir8: in std_logic;
      ir10: in std_logic;
      ir11: in std_logic;
      ir19: in std_logic;
      ir20: in std_logic;
      ir21: in std_logic;
      ir22: in std_logic;
      ir23: in std_logic;
      ir25: in std_logic;
      ir26: in std_logic;
      ir27: in std_logic;
      ir28: in std_logic;
      ir29: in std_logic;
      ir43: in std_logic;
      ir44: in std_logic;
      \-ir31\: in std_logic;
      nop: in std_logic;
      dest: out std_logic;
      \-destimod0\: out std_logic;
      \-destimod1\: out std_logic;
      \-destintctl\: out std_logic;
      \-destlc\: out std_logic;
      destm: out std_logic;
      \-destmdr\: out std_logic;
      \-destmem\: out std_logic;
      \-destpdl(p)\: out std_logic;
      \-destpdl(x)\: out std_logic;
      \-destpdlp\: out std_logic;
      \-destpdltop\: out std_logic;
      \-destpdlx\: out std_logic;
      \-destspc\: out std_logic;
      \-destvma\: out std_logic;
      \-div\: out std_logic;
      \-funct2\: out std_logic;
      imod: out std_logic;
      \-iralu\: out std_logic;
      \-irbyte\: out std_logic;
      irdisp: out std_logic;
      \-irdisp\: out std_logic;
      irjump: out std_logic;
      \-irjump\: out std_logic;
      \-mul\: out std_logic;
      \-srcdc\: out std_logic;
      \-srclc\: out std_logic;
      \-srcmap\: out std_logic;
      \-srcmd\: out std_logic;
      \-srcopc\: out std_logic;
      \-srcpdlidx\: out std_logic;
      \-srcpdlpop\: out std_logic;
      \-srcpdlptr\: out std_logic;
      \-srcpdltop\: out std_logic;
      \-srcq\: out std_logic;
      \-srcspc\: out std_logic;
      \-srcspcpop\: out std_logic;
      \-srcvma\: out std_logic
    );
  end component;
  component dmem_set is
      -- internal signals: aa16 aa17 dadr10a dadr10c \-dadr10a\ 
      -- internal signals: \-dadr10c\ dispwr \-dmapbenb\ dmask0 dmask1 
      -- internal signals: dmask2 dmask3 dmask4 dmask5 dmask6 
      -- internal signals: dpar ir8b ir9b ir12b ir13b 
      -- internal signals: ir14b ir15b ir16b ir17b ir18b 
      -- internal signals: ir19b ir20b ir21b ir22b vmo18 
      -- internal signals: vmo19 
    port (
      a0: in std_logic;
      a1: in std_logic;
      a2: in std_logic;
      a3: in std_logic;
      a4: in std_logic;
      a5: in std_logic;
      a6: in std_logic;
      a7: in std_logic;
      a8: in std_logic;
      a9: in std_logic;
      a10: in std_logic;
      a11: in std_logic;
      a12: in std_logic;
      a13: in std_logic;
      a14: in std_logic;
      a15: in std_logic;
      a16: in std_logic;
      a17: in std_logic;
      clk3e: in std_logic;
      dispenb: in std_logic;
      \-funct2\: in std_logic;
      hi4: in std_logic;
      hi6: in std_logic;
      hi11: in std_logic;
      ir5: in std_logic;
      ir6: in std_logic;
      ir7: in std_logic;
      ir8: in std_logic;
      ir9: in std_logic;
      ir12: in std_logic;
      ir13: in std_logic;
      ir14: in std_logic;
      ir15: in std_logic;
      ir16: in std_logic;
      ir17: in std_logic;
      ir18: in std_logic;
      ir19: in std_logic;
      ir20: in std_logic;
      ir21: in std_logic;
      ir22: in std_logic;
      ir32: in std_logic;
      ir33: in std_logic;
      ir34: in std_logic;
      ir35: in std_logic;
      ir36: in std_logic;
      ir37: in std_logic;
      ir38: in std_logic;
      ir39: in std_logic;
      ir40: in std_logic;
      ir41: in std_logic;
      \-irdisp\: in std_logic;
      r0: in std_logic;
      r1: in std_logic;
      r2: in std_logic;
      r3: in std_logic;
      r4: in std_logic;
      r5: in std_logic;
      r6: in std_logic;
      wp2: in std_logic;
      dn: inout std_logic;
      dpc0: inout std_logic;
      dpc1: inout std_logic;
      dpc2: inout std_logic;
      dpc3: inout std_logic;
      dpc5: inout std_logic;
      dpc6: inout std_logic;
      dpc7: inout std_logic;
      dpc8: inout std_logic;
      dpc9: inout std_logic;
      dpc10: inout std_logic;
      dpc11: inout std_logic;
      dpc12: inout std_logic;
      dpc13: inout std_logic;
      aa0: out std_logic;
      aa1: out std_logic;
      aa2: out std_logic;
      aa3: out std_logic;
      aa4: out std_logic;
      aa5: out std_logic;
      aa6: out std_logic;
      aa7: out std_logic;
      aa8: out std_logic;
      aa9: out std_logic;
      aa10: out std_logic;
      aa11: out std_logic;
      aa12: out std_logic;
      aa13: out std_logic;
      aa14: out std_logic;
      aa15: out std_logic;
      dc0: out std_logic;
      dc1: out std_logic;
      dc2: out std_logic;
      dc3: out std_logic;
      dc4: out std_logic;
      dc5: out std_logic;
      dc6: out std_logic;
      dc7: out std_logic;
      dc8: out std_logic;
      dc9: out std_logic;
      dp: out std_logic;
      dparok: out std_logic;
      dpc4: out std_logic;
      dr: out std_logic;
      \-vmo18\: out std_logic;
      \-vmo19\: out std_logic
    );
  end component;
  component fetch_set is

    port (
      aa0: in std_logic;
      aa1: in std_logic;
      aa2: in std_logic;
      aa3: in std_logic;
      aa4: in std_logic;
      aa5: in std_logic;
      aa6: in std_logic;
      aa7: in std_logic;
      aa8: in std_logic;
      aa9: in std_logic;
      aa10: in std_logic;
      aa11: in std_logic;
      aa12: in std_logic;
      aa13: in std_logic;
      aa14: in std_logic;
      aa15: in std_logic;
      clk2c: in std_logic;
      clk4c: in std_logic;
      \-idebug\: in std_logic;
      \-lddbirh\: in std_logic;
      \-lddbirl\: in std_logic;
      \-lddbirm\: in std_logic;
      m0: in std_logic;
      m1: in std_logic;
      m2: in std_logic;
      m3: in std_logic;
      m4: in std_logic;
      m5: in std_logic;
      m6: in std_logic;
      m7: in std_logic;
      m8: in std_logic;
      m9: in std_logic;
      m10: in std_logic;
      m11: in std_logic;
      m12: in std_logic;
      m13: in std_logic;
      m14: in std_logic;
      m15: in std_logic;
      m16: in std_logic;
      m17: in std_logic;
      m18: in std_logic;
      m19: in std_logic;
      m20: in std_logic;
      m21: in std_logic;
      m22: in std_logic;
      m23: in std_logic;
      m24: in std_logic;
      m25: in std_logic;
      m26: in std_logic;
      m27: in std_logic;
      m28: in std_logic;
      m29: in std_logic;
      m30: in std_logic;
      m31: in std_logic;
      spy0: in std_logic;
      spy1: in std_logic;
      spy2: in std_logic;
      spy3: in std_logic;
      spy4: in std_logic;
      spy5: in std_logic;
      spy6: in std_logic;
      spy7: in std_logic;
      spy8: in std_logic;
      spy9: in std_logic;
      spy10: in std_logic;
      spy11: in std_logic;
      spy12: in std_logic;
      spy13: in std_logic;
      spy14: in std_logic;
      spy15: in std_logic;
      i0: out std_logic;
      i1: out std_logic;
      i2: out std_logic;
      i3: out std_logic;
      i4: out std_logic;
      i5: out std_logic;
      i6: out std_logic;
      i7: out std_logic;
      i8: out std_logic;
      i9: out std_logic;
      i10: out std_logic;
      i11: out std_logic;
      i12: out std_logic;
      i13: out std_logic;
      i14: out std_logic;
      i15: out std_logic;
      i16: out std_logic;
      i17: out std_logic;
      i18: out std_logic;
      i19: out std_logic;
      i20: out std_logic;
      i21: out std_logic;
      i22: out std_logic;
      i23: out std_logic;
      i24: out std_logic;
      i25: out std_logic;
      i26: out std_logic;
      i27: out std_logic;
      i28: out std_logic;
      i29: out std_logic;
      i30: out std_logic;
      i31: out std_logic;
      i32: out std_logic;
      i33: out std_logic;
      i34: out std_logic;
      i35: out std_logic;
      i36: out std_logic;
      i37: out std_logic;
      i38: out std_logic;
      i39: out std_logic;
      i40: out std_logic;
      i41: out std_logic;
      i42: out std_logic;
      i43: out std_logic;
      i44: out std_logic;
      i45: out std_logic;
      i46: out std_logic;
      i47: out std_logic;
      iwr0: out std_logic;
      iwr1: out std_logic;
      iwr2: out std_logic;
      iwr3: out std_logic;
      iwr4: out std_logic;
      iwr5: out std_logic;
      iwr6: out std_logic;
      iwr7: out std_logic;
      iwr8: out std_logic;
      iwr9: out std_logic;
      iwr10: out std_logic;
      iwr11: out std_logic;
      iwr12: out std_logic;
      iwr13: out std_logic;
      iwr14: out std_logic;
      iwr15: out std_logic;
      iwr16: out std_logic;
      iwr17: out std_logic;
      iwr18: out std_logic;
      iwr19: out std_logic;
      iwr20: out std_logic;
      iwr21: out std_logic;
      iwr22: out std_logic;
      iwr23: out std_logic;
      iwr24: out std_logic;
      iwr25: out std_logic;
      iwr26: out std_logic;
      iwr27: out std_logic;
      iwr28: out std_logic;
      iwr29: out std_logic;
      iwr30: out std_logic;
      iwr31: out std_logic;
      iwr32: out std_logic;
      iwr33: out std_logic;
      iwr34: out std_logic;
      iwr35: out std_logic;
      iwr36: out std_logic;
      iwr37: out std_logic;
      iwr38: out std_logic;
      iwr39: out std_logic;
      iwr40: out std_logic;
      iwr41: out std_logic;
      iwr42: out std_logic;
      iwr43: out std_logic;
      iwr44: out std_logic;
      iwr45: out std_logic;
      iwr46: out std_logic;
      iwr47: out std_logic;
      iwr48: out std_logic
    );
  end component;
  component flowc_set is

    port (
      clk3c: in std_logic;
      dp: in std_logic;
      dr: in std_logic;
      \-funct2\: in std_logic;
      hi4: in std_logic;
      ir6: in std_logic;
      ir7: in std_logic;
      ir8: in std_logic;
      ir9: in std_logic;
      ir42: in std_logic;
      irdisp: in std_logic;
      \-irdisp\: in std_logic;
      irjump: in std_logic;
      jcond: in std_logic;
      \-jcond\: in std_logic;
      \-nop11\: in std_logic;
      \-reset\: in std_logic;
      \-srcspc\: in std_logic;
      \-srcspcpop\: in std_logic;
      \-trap\: in std_logic;
      tse3a: in std_logic;
      wp4c: in std_logic;
      \-destspc\: out std_logic;
      destspcd: out std_logic;
      dispenb: out std_logic;
      dn: out std_logic;
      iwrited: out std_logic;
      \-iwrited\: out std_logic;
      n: out std_logic;
      nop: out std_logic;
      \-nopa\: out std_logic;
      pcs0: out std_logic;
      pcs1: out std_logic;
      spcdrive: out std_logic;
      \-spcdrive\: out std_logic;
      spcenb: out std_logic;
      \-spcnt\: out std_logic;
      \-spcpass\: out std_logic;
      spcwpass: out std_logic;
      \-spcwpass\: out std_logic;
      \-spop\: out std_logic;
      spush: out std_logic;
      spushd: out std_logic;
      \-srcspcpopreal\: out std_logic;
      \-swpa\: out std_logic;
      \-swpb\: out std_logic
    );
  end component;
  component imem_set is
      -- internal signals: \-ice0a\ \-ice0b\ \-ice0c\ \-ice0d\ \-ice1a\ 
      -- internal signals: \-ice1b\ \-ice1c\ \-ice1d\ \-ice2a\ \-ice2b\ 
      -- internal signals: \-ice2c\ \-ice2d\ \-ice3a\ \-ice3b\ \-ice3c\ 
      -- internal signals: \-ice3d\ \-iwea\ \-iweb\ \-iwec\ \-iwed\ 
      -- internal signals: \-iwee\ \-iwef\ \-iweg\ \-iweh\ \-iwei\ 
      -- internal signals: \-iwej\ \-iwek\ \-iwel\ \-iwem\ \-iwen\ 
      -- internal signals: \-iweo\ \-iwep\ \-pcb0\ \-pcb1\ \-pcb2\ 
      -- internal signals: \-pcb3\ \-pcb4\ \-pcb5\ \-pcb6\ \-pcb7\ 
      -- internal signals: \-pcb8\ \-pcb9\ \-pcb10\ \-pcb11\ \-pcc0\ 
      -- internal signals: \-pcc1\ \-pcc2\ \-pcc3\ \-pcc4\ \-pcc5\ 
      -- internal signals: \-pcc6\ \-pcc7\ \-pcc8\ \-pcc9\ \-pcc10\ 
      -- internal signals: \-pcc11\ 
    port (
      hi1: in std_logic;
      idebug: in std_logic;
      iwr0: in std_logic;
      iwr1: in std_logic;
      iwr2: in std_logic;
      iwr3: in std_logic;
      iwr4: in std_logic;
      iwr5: in std_logic;
      iwr6: in std_logic;
      iwr7: in std_logic;
      iwr8: in std_logic;
      iwr9: in std_logic;
      iwr10: in std_logic;
      iwr11: in std_logic;
      iwr12: in std_logic;
      iwr13: in std_logic;
      iwr14: in std_logic;
      iwr15: in std_logic;
      iwr16: in std_logic;
      iwr17: in std_logic;
      iwr18: in std_logic;
      iwr19: in std_logic;
      iwr20: in std_logic;
      iwr21: in std_logic;
      iwr22: in std_logic;
      iwr23: in std_logic;
      iwr24: in std_logic;
      iwr25: in std_logic;
      iwr26: in std_logic;
      iwr27: in std_logic;
      iwr28: in std_logic;
      iwr29: in std_logic;
      iwr30: in std_logic;
      iwr31: in std_logic;
      iwr32: in std_logic;
      iwr33: in std_logic;
      iwr34: in std_logic;
      iwr35: in std_logic;
      iwr36: in std_logic;
      iwr37: in std_logic;
      iwr38: in std_logic;
      iwr39: in std_logic;
      iwr40: in std_logic;
      iwr41: in std_logic;
      iwr42: in std_logic;
      iwr43: in std_logic;
      iwr44: in std_logic;
      iwr45: in std_logic;
      iwr46: in std_logic;
      iwr47: in std_logic;
      iwr48: in std_logic;
      \-iwrited\: in std_logic;
      pc0: in std_logic;
      pc1: in std_logic;
      pc2: in std_logic;
      pc3: in std_logic;
      pc4: in std_logic;
      pc5: in std_logic;
      pc6: in std_logic;
      pc7: in std_logic;
      pc8: in std_logic;
      pc9: in std_logic;
      pc10: in std_logic;
      pc11: in std_logic;
      pc12: in std_logic;
      pc13: in std_logic;
      promdisabled: in std_logic;
      \-wp5\: in std_logic;
      i0: out std_logic;
      i1: out std_logic;
      i2: out std_logic;
      i3: out std_logic;
      i4: out std_logic;
      i5: out std_logic;
      i6: out std_logic;
      i7: out std_logic;
      i8: out std_logic;
      i9: out std_logic;
      i10: out std_logic;
      i11: out std_logic;
      i12: out std_logic;
      i13: out std_logic;
      i14: out std_logic;
      i15: out std_logic;
      i16: out std_logic;
      i17: out std_logic;
      i18: out std_logic;
      i19: out std_logic;
      i20: out std_logic;
      i21: out std_logic;
      i22: out std_logic;
      i23: out std_logic;
      i24: out std_logic;
      i25: out std_logic;
      i26: out std_logic;
      i27: out std_logic;
      i28: out std_logic;
      i29: out std_logic;
      i30: out std_logic;
      i31: out std_logic;
      i32: out std_logic;
      i33: out std_logic;
      i34: out std_logic;
      i35: out std_logic;
      i36: out std_logic;
      i37: out std_logic;
      i38: out std_logic;
      i39: out std_logic;
      i40: out std_logic;
      i41: out std_logic;
      i42: out std_logic;
      i43: out std_logic;
      i44: out std_logic;
      i45: out std_logic;
      i46: out std_logic;
      i47: out std_logic;
      i48: out std_logic;
      \-iwriteda\: out std_logic;
      \-promdisabled\: out std_logic
    );
  end component;
  component ireg_set is
      -- internal signals: iob0 iob1 iob2 iob3 iob4 
      -- internal signals: iob5 iob6 iob7 iob8 iob9 
      -- internal signals: iob10 iob11 iob12 iob13 iob14 
      -- internal signals: iob15 iob16 iob17 iob18 iob19 
      -- internal signals: iob20 iob21 iob22 iob23 iob24 
      -- internal signals: iob25 iob26 iob27 iob28 iob29 
      -- internal signals: iob30 iob31 iob32 iob33 iob34 
      -- internal signals: iob35 iob36 iob37 iob38 iob39 
      -- internal signals: iob40 iob41 iob42 iob43 iob44 
      -- internal signals: iob45 iob46 iob47 
    port (
      clk3a: in std_logic;
      clk3b: in std_logic;
      \-destimod0\: in std_logic;
      \-destimod1\: in std_logic;
      i0: in std_logic;
      i1: in std_logic;
      i2: in std_logic;
      i3: in std_logic;
      i4: in std_logic;
      i5: in std_logic;
      i6: in std_logic;
      i7: in std_logic;
      i8: in std_logic;
      i9: in std_logic;
      i10: in std_logic;
      i11: in std_logic;
      i12: in std_logic;
      i13: in std_logic;
      i14: in std_logic;
      i15: in std_logic;
      i16: in std_logic;
      i17: in std_logic;
      i18: in std_logic;
      i19: in std_logic;
      i20: in std_logic;
      i21: in std_logic;
      i22: in std_logic;
      i23: in std_logic;
      i24: in std_logic;
      i25: in std_logic;
      i26: in std_logic;
      i27: in std_logic;
      i28: in std_logic;
      i29: in std_logic;
      i30: in std_logic;
      i31: in std_logic;
      i32: in std_logic;
      i33: in std_logic;
      i34: in std_logic;
      i35: in std_logic;
      i36: in std_logic;
      i37: in std_logic;
      i38: in std_logic;
      i39: in std_logic;
      i40: in std_logic;
      i41: in std_logic;
      i42: in std_logic;
      i43: in std_logic;
      i44: in std_logic;
      i45: in std_logic;
      i46: in std_logic;
      i47: in std_logic;
      i48: in std_logic;
      imodd: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      ob10: in std_logic;
      ob11: in std_logic;
      ob12: in std_logic;
      ob13: in std_logic;
      ob14: in std_logic;
      ob15: in std_logic;
      ob16: in std_logic;
      ob17: in std_logic;
      ob18: in std_logic;
      ob19: in std_logic;
      ob20: in std_logic;
      ob21: in std_logic;
      ob22: in std_logic;
      ob23: in std_logic;
      ob24: in std_logic;
      ob25: in std_logic;
      iparok: out std_logic;
      ir0: out std_logic;
      ir1: out std_logic;
      ir2: out std_logic;
      ir3: out std_logic;
      ir4: out std_logic;
      ir5: out std_logic;
      ir6: out std_logic;
      ir7: out std_logic;
      ir8: out std_logic;
      ir9: out std_logic;
      ir10: out std_logic;
      ir11: out std_logic;
      ir12: out std_logic;
      ir13: out std_logic;
      ir14: out std_logic;
      ir15: out std_logic;
      ir16: out std_logic;
      ir17: out std_logic;
      ir18: out std_logic;
      ir19: out std_logic;
      ir20: out std_logic;
      ir21: out std_logic;
      ir22: out std_logic;
      ir23: out std_logic;
      ir24: out std_logic;
      ir25: out std_logic;
      ir26: out std_logic;
      ir27: out std_logic;
      ir28: out std_logic;
      ir29: out std_logic;
      ir30: out std_logic;
      ir31: out std_logic;
      ir32: out std_logic;
      ir33: out std_logic;
      ir34: out std_logic;
      ir35: out std_logic;
      ir36: out std_logic;
      ir37: out std_logic;
      ir38: out std_logic;
      ir39: out std_logic;
      ir40: out std_logic;
      ir41: out std_logic;
      ir42: out std_logic;
      ir43: out std_logic;
      ir44: out std_logic;
      ir45: out std_logic;
      ir46: out std_logic;
      ir47: out std_logic;
      ir48: out std_logic
    );
  end component;
  component jumpc_set is

    port (
      \a=m\: in std_logic;
      alu32: in std_logic;
      clk3c: in std_logic;
      \-destintctl\: in std_logic;
      hi4: in std_logic;
      ir0: in std_logic;
      ir1: in std_logic;
      ir2: in std_logic;
      ir5: in std_logic;
      ir45: in std_logic;
      ir46: in std_logic;
      \-nopa\: in std_logic;
      ob26: in std_logic;
      ob27: in std_logic;
      ob28: in std_logic;
      ob29: in std_logic;
      r0: in std_logic;
      \-reset\: in std_logic;
      sintr: in std_logic;
      \-vmaok\: in std_logic;
      \-ilong\: out std_logic;
      \int.enable\: out std_logic;
      jcond: out std_logic;
      \-jcond\: out std_logic;
      \lc byte mode\: out std_logic;
      \prog.unibus.reset\: out std_logic;
      \sequence.break\: out std_logic;
      \-statbit\: out std_logic
    );
  end component;
  component lcreg_set is
      -- internal signals: lc1 lc0b 
    port (
      clk1a: in std_logic;
      clk2a: in std_logic;
      clk2c: in std_logic;
      clk3c: in std_logic;
      \-destlc\: in std_logic;
      hi11: in std_logic;
      \int.enable\: in std_logic;
      ir10: in std_logic;
      ir11: in std_logic;
      ir24: in std_logic;
      \-ir3\: in std_logic;
      \-ir4\: in std_logic;
      irdisp: in std_logic;
      \lc byte mode\: in std_logic;
      \-lcry3\: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      ob10: in std_logic;
      ob11: in std_logic;
      ob12: in std_logic;
      ob13: in std_logic;
      ob14: in std_logic;
      ob15: in std_logic;
      ob16: in std_logic;
      ob17: in std_logic;
      ob18: in std_logic;
      ob19: in std_logic;
      ob20: in std_logic;
      ob21: in std_logic;
      ob22: in std_logic;
      ob23: in std_logic;
      ob24: in std_logic;
      ob25: in std_logic;
      \prog.unibus.reset\: in std_logic;
      \-reset\: in std_logic;
      \sequence.break\: in std_logic;
      spc1: in std_logic;
      spc14: in std_logic;
      \-spop\: in std_logic;
      \-srclc\: in std_logic;
      \-srcspcpopreal\: in std_logic;
      tse1a: in std_logic;
      \-ifetch\: out std_logic;
      lc2: out std_logic;
      lc3: out std_logic;
      lc4: out std_logic;
      lc5: out std_logic;
      lc6: out std_logic;
      lc7: out std_logic;
      lc8: out std_logic;
      lc9: out std_logic;
      lc10: out std_logic;
      lc11: out std_logic;
      lc12: out std_logic;
      lc13: out std_logic;
      lc14: out std_logic;
      lc15: out std_logic;
      lc16: out std_logic;
      lc17: out std_logic;
      lc18: out std_logic;
      lc19: out std_logic;
      lc20: out std_logic;
      lc21: out std_logic;
      lc22: out std_logic;
      lc23: out std_logic;
      lc24: out std_logic;
      lc25: out std_logic;
      lcinc: out std_logic;
      lcry3: out std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mf12: out std_logic;
      mf13: out std_logic;
      mf14: out std_logic;
      mf15: out std_logic;
      mf16: out std_logic;
      mf17: out std_logic;
      mf18: out std_logic;
      mf19: out std_logic;
      mf20: out std_logic;
      mf21: out std_logic;
      mf22: out std_logic;
      mf23: out std_logic;
      mf24: out std_logic;
      mf25: out std_logic;
      mf26: out std_logic;
      mf27: out std_logic;
      mf28: out std_logic;
      mf29: out std_logic;
      mf30: out std_logic;
      mf31: out std_logic;
      needfetch: out std_logic;
      \-sh3\: out std_logic;
      \-sh4\: out std_logic;
      sintr: out std_logic;
      spc1a: out std_logic
    );
  end component;
  component lreg_set is

    port (
      clk3f: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      ob10: in std_logic;
      ob11: in std_logic;
      ob12: in std_logic;
      ob13: in std_logic;
      ob14: in std_logic;
      ob15: in std_logic;
      ob16: in std_logic;
      ob17: in std_logic;
      ob18: in std_logic;
      ob19: in std_logic;
      ob20: in std_logic;
      ob21: in std_logic;
      ob22: in std_logic;
      ob23: in std_logic;
      ob24: in std_logic;
      ob25: in std_logic;
      ob26: in std_logic;
      ob27: in std_logic;
      ob28: in std_logic;
      ob29: in std_logic;
      ob30: in std_logic;
      ob31: in std_logic;
      l0: out std_logic;
      l1: out std_logic;
      l2: out std_logic;
      l3: out std_logic;
      l4: out std_logic;
      l5: out std_logic;
      l6: out std_logic;
      l7: out std_logic;
      l8: out std_logic;
      l9: out std_logic;
      l10: out std_logic;
      l11: out std_logic;
      l12: out std_logic;
      l13: out std_logic;
      l14: out std_logic;
      l15: out std_logic;
      l16: out std_logic;
      l17: out std_logic;
      l18: out std_logic;
      l19: out std_logic;
      l20: out std_logic;
      l21: out std_logic;
      l22: out std_logic;
      l23: out std_logic;
      l24: out std_logic;
      l25: out std_logic;
      l26: out std_logic;
      l27: out std_logic;
      l28: out std_logic;
      l29: out std_logic;
      l30: out std_logic;
      l31: out std_logic;
      lparity: out std_logic
    );
  end component;
  component md_set is
      -- internal signals: \-mds0\ \-mds1\ \-mds2\ \-mds3\ \-mds4\ 
      -- internal signals: \-mds5\ \-mds6\ \-mds7\ \-mds8\ \-mds9\ 
      -- internal signals: \-mds10\ \-mds11\ \-mds12\ \-mds13\ \-mds14\ 
      -- internal signals: \-mds15\ \-mds16\ \-mds17\ \-mds18\ \-mds19\ 
      -- internal signals: \-mds20\ \-mds21\ \-mds22\ \-mds23\ \-mds24\ 
      -- internal signals: \-mds25\ \-mds26\ \-mds27\ \-mds28\ \-mds29\ 
      -- internal signals: \-mds30\ \-mds31\ 
    port (
      \-clk2c\: in std_logic;
      \-destmdr\: in std_logic;
      hi11: in std_logic;
      mdparodd: in std_logic;
      mdsela: in std_logic;
      mdselb: in std_logic;
      \-memdrive.a\: in std_logic;
      \-memdrive.b\: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      ob10: in std_logic;
      ob11: in std_logic;
      ob12: in std_logic;
      ob13: in std_logic;
      ob14: in std_logic;
      ob15: in std_logic;
      ob16: in std_logic;
      ob17: in std_logic;
      ob18: in std_logic;
      ob19: in std_logic;
      ob20: in std_logic;
      ob21: in std_logic;
      ob22: in std_logic;
      ob23: in std_logic;
      ob24: in std_logic;
      ob25: in std_logic;
      ob26: in std_logic;
      ob27: in std_logic;
      ob28: in std_logic;
      ob29: in std_logic;
      ob30: in std_logic;
      ob31: in std_logic;
      \-srcmd\: in std_logic;
      tse2: in std_logic;
      \-md0\: out std_logic;
      \-md1\: out std_logic;
      \-md2\: out std_logic;
      \-md3\: out std_logic;
      \-md4\: out std_logic;
      \-md5\: out std_logic;
      \-md6\: out std_logic;
      \-md7\: out std_logic;
      \-md8\: out std_logic;
      \-md9\: out std_logic;
      \-md10\: out std_logic;
      \-md11\: out std_logic;
      \-md12\: out std_logic;
      \-md13\: out std_logic;
      \-md14\: out std_logic;
      \-md15\: out std_logic;
      \-md16\: out std_logic;
      \-md17\: out std_logic;
      \-md18\: out std_logic;
      \-md19\: out std_logic;
      \-md20\: out std_logic;
      \-md21\: out std_logic;
      \-md22\: out std_logic;
      \-md23\: out std_logic;
      \-md24\: out std_logic;
      \-md25\: out std_logic;
      \-md26\: out std_logic;
      \-md27\: out std_logic;
      \-md28\: out std_logic;
      \-md29\: out std_logic;
      \-md30\: out std_logic;
      \-md31\: out std_logic;
      mdhaspar: out std_logic;
      mdpar: out std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mf12: out std_logic;
      mf13: out std_logic;
      mf14: out std_logic;
      mf15: out std_logic;
      mf16: out std_logic;
      mf17: out std_logic;
      mf18: out std_logic;
      mf19: out std_logic;
      mf20: out std_logic;
      mf21: out std_logic;
      mf22: out std_logic;
      mf23: out std_logic;
      mf24: out std_logic;
      mf25: out std_logic;
      mf26: out std_logic;
      mf27: out std_logic;
      mf28: out std_logic;
      mf29: out std_logic;
      mf30: out std_logic;
      mf31: out std_logic
    );
  end component;
  component mmem_set is
      -- internal signals: \-madr0a\ \-madr0b\ \-madr1a\ \-madr1b\ \-madr2a\ 
      -- internal signals: \-madr2b\ \-madr3a\ \-madr3b\ \-madr4a\ \-madr4b\ 
      -- internal signals: mmem2 mmem3 mmem5 mmem7 mmem9 
      -- internal signals: mmem11 mmem13 mmem15 mmem17 mmem19 
      -- internal signals: mmem21 mmem23 mmem25 mmem27 mmem29 
      -- internal signals: mmem31 \-mpass\ mpassl \-mpassl\ \-mpassm\ 
      -- internal signals: \-mwpa\ \-mwpb\ 
    port (
      clk4a: in std_logic;
      clk4e: in std_logic;
      destmd: in std_logic;
      hi2: in std_logic;
      hi3: in std_logic;
      ir26: in std_logic;
      ir27: in std_logic;
      ir28: in std_logic;
      ir29: in std_logic;
      ir30: in std_logic;
      \-ir31\: in std_logic;
      l0: in std_logic;
      l1: in std_logic;
      l2: in std_logic;
      l3: in std_logic;
      l4: in std_logic;
      l5: in std_logic;
      l6: in std_logic;
      l7: in std_logic;
      l8: in std_logic;
      l9: in std_logic;
      l10: in std_logic;
      l11: in std_logic;
      l12: in std_logic;
      l13: in std_logic;
      l14: in std_logic;
      l15: in std_logic;
      l16: in std_logic;
      l17: in std_logic;
      l18: in std_logic;
      l19: in std_logic;
      l20: in std_logic;
      l21: in std_logic;
      l22: in std_logic;
      l23: in std_logic;
      l24: in std_logic;
      l25: in std_logic;
      l26: in std_logic;
      l27: in std_logic;
      l28: in std_logic;
      l29: in std_logic;
      l30: in std_logic;
      l31: in std_logic;
      lparity: in std_logic;
      pdlenb: in std_logic;
      spcenb: in std_logic;
      tse1a: in std_logic;
      tse4a: in std_logic;
      wadr0: in std_logic;
      wadr1: in std_logic;
      wadr2: in std_logic;
      wadr3: in std_logic;
      wadr4: in std_logic;
      wp4b: in std_logic;
      mf0: inout std_logic;
      mf1: inout std_logic;
      mf2: inout std_logic;
      mf3: inout std_logic;
      mf4: inout std_logic;
      mf5: inout std_logic;
      mf6: inout std_logic;
      mf7: inout std_logic;
      mf8: inout std_logic;
      mf9: inout std_logic;
      mf10: inout std_logic;
      mf11: inout std_logic;
      mf12: inout std_logic;
      mf13: inout std_logic;
      mf14: inout std_logic;
      mf15: inout std_logic;
      mf16: inout std_logic;
      mf17: inout std_logic;
      mf18: inout std_logic;
      mf19: inout std_logic;
      mf20: inout std_logic;
      mf21: inout std_logic;
      mf22: inout std_logic;
      mf23: inout std_logic;
      mf24: inout std_logic;
      mf25: inout std_logic;
      mf26: inout std_logic;
      mf27: inout std_logic;
      mf28: inout std_logic;
      mf29: inout std_logic;
      mf30: inout std_logic;
      mf31: inout std_logic;
      m0: out std_logic;
      m1: out std_logic;
      m2: out std_logic;
      m3: out std_logic;
      m4: out std_logic;
      m5: out std_logic;
      m6: out std_logic;
      m7: out std_logic;
      m8: out std_logic;
      m9: out std_logic;
      m10: out std_logic;
      m11: out std_logic;
      m12: out std_logic;
      m13: out std_logic;
      m14: out std_logic;
      m15: out std_logic;
      m16: out std_logic;
      m17: out std_logic;
      m18: out std_logic;
      m19: out std_logic;
      m20: out std_logic;
      m21: out std_logic;
      m22: out std_logic;
      m23: out std_logic;
      m24: out std_logic;
      m25: out std_logic;
      m26: out std_logic;
      m27: out std_logic;
      m28: out std_logic;
      m29: out std_logic;
      m30: out std_logic;
      m31: out std_logic;
      mparity: out std_logic;
      srcm: out std_logic
    );
  end component;
  component mos_set is

    port (
      a0: in std_logic;
      a1: in std_logic;
      a2: in std_logic;
      a3: in std_logic;
      a4: in std_logic;
      a5: in std_logic;
      a6: in std_logic;
      a7: in std_logic;
      a8: in std_logic;
      a9: in std_logic;
      a10: in std_logic;
      a11: in std_logic;
      a12: in std_logic;
      a13: in std_logic;
      a14: in std_logic;
      a15: in std_logic;
      a16: in std_logic;
      a17: in std_logic;
      a18: in std_logic;
      a19: in std_logic;
      a20: in std_logic;
      a21: in std_logic;
      a22: in std_logic;
      a23: in std_logic;
      a24: in std_logic;
      a25: in std_logic;
      a26: in std_logic;
      a27: in std_logic;
      a28: in std_logic;
      a29: in std_logic;
      a30: in std_logic;
      a31b: in std_logic;
      alu0: in std_logic;
      alu1: in std_logic;
      alu2: in std_logic;
      alu3: in std_logic;
      alu4: in std_logic;
      alu5: in std_logic;
      alu6: in std_logic;
      alu7: in std_logic;
      alu8: in std_logic;
      alu9: in std_logic;
      alu10: in std_logic;
      alu11: in std_logic;
      alu12: in std_logic;
      alu13: in std_logic;
      alu14: in std_logic;
      alu15: in std_logic;
      alu16: in std_logic;
      alu17: in std_logic;
      alu18: in std_logic;
      alu19: in std_logic;
      alu20: in std_logic;
      alu21: in std_logic;
      alu22: in std_logic;
      alu23: in std_logic;
      alu24: in std_logic;
      alu25: in std_logic;
      alu26: in std_logic;
      alu27: in std_logic;
      alu28: in std_logic;
      alu29: in std_logic;
      alu30: in std_logic;
      alu31: in std_logic;
      alu32: in std_logic;
      msk0: in std_logic;
      msk1: in std_logic;
      msk2: in std_logic;
      msk3: in std_logic;
      msk4: in std_logic;
      msk5: in std_logic;
      msk6: in std_logic;
      msk7: in std_logic;
      msk8: in std_logic;
      msk9: in std_logic;
      msk10: in std_logic;
      msk11: in std_logic;
      msk12: in std_logic;
      msk13: in std_logic;
      msk14: in std_logic;
      msk15: in std_logic;
      msk16: in std_logic;
      msk17: in std_logic;
      msk18: in std_logic;
      msk19: in std_logic;
      msk20: in std_logic;
      msk21: in std_logic;
      msk22: in std_logic;
      msk23: in std_logic;
      msk24: in std_logic;
      msk25: in std_logic;
      msk26: in std_logic;
      msk27: in std_logic;
      msk28: in std_logic;
      msk29: in std_logic;
      msk30: in std_logic;
      msk31: in std_logic;
      osel0a: in std_logic;
      osel0b: in std_logic;
      osel1a: in std_logic;
      osel1b: in std_logic;
      q31: in std_logic;
      r0: in std_logic;
      r1: in std_logic;
      r2: in std_logic;
      r3: in std_logic;
      r4: in std_logic;
      r5: in std_logic;
      r6: in std_logic;
      r7: in std_logic;
      r8: in std_logic;
      r9: in std_logic;
      r10: in std_logic;
      r11: in std_logic;
      r12: in std_logic;
      r13: in std_logic;
      r14: in std_logic;
      r15: in std_logic;
      r16: in std_logic;
      r17: in std_logic;
      r18: in std_logic;
      r19: in std_logic;
      r20: in std_logic;
      r21: in std_logic;
      r22: in std_logic;
      r23: in std_logic;
      r24: in std_logic;
      r25: in std_logic;
      r26: in std_logic;
      r27: in std_logic;
      r28: in std_logic;
      r29: in std_logic;
      r30: in std_logic;
      r31: in std_logic;
      ob0: out std_logic;
      ob1: out std_logic;
      ob2: out std_logic;
      ob3: out std_logic;
      ob4: out std_logic;
      ob5: out std_logic;
      ob6: out std_logic;
      ob7: out std_logic;
      ob8: out std_logic;
      ob9: out std_logic;
      ob10: out std_logic;
      ob11: out std_logic;
      ob12: out std_logic;
      ob13: out std_logic;
      ob14: out std_logic;
      ob15: out std_logic;
      ob16: out std_logic;
      ob17: out std_logic;
      ob18: out std_logic;
      ob19: out std_logic;
      ob20: out std_logic;
      ob21: out std_logic;
      ob22: out std_logic;
      ob23: out std_logic;
      ob24: out std_logic;
      ob25: out std_logic;
      ob26: out std_logic;
      ob27: out std_logic;
      ob28: out std_logic;
      ob29: out std_logic;
      ob30: out std_logic;
      ob31: out std_logic
    );
  end component;
  component npc_set is

    port (
      clk4b: in std_logic;
      dpc4: in std_logic;
      hi4: in std_logic;
      ir12: in std_logic;
      ir13: in std_logic;
      ir14: in std_logic;
      ir15: in std_logic;
      ir16: in std_logic;
      ir17: in std_logic;
      ir18: in std_logic;
      ir19: in std_logic;
      ir20: in std_logic;
      ir21: in std_logic;
      ir22: in std_logic;
      ir23: in std_logic;
      ir24: in std_logic;
      ir25: in std_logic;
      pcs0: in std_logic;
      pcs1: in std_logic;
      spc1a: in std_logic;
      trapa: in std_logic;
      trapb: in std_logic;
      dpc0: out std_logic;
      dpc1: out std_logic;
      dpc2: out std_logic;
      dpc3: out std_logic;
      dpc5: out std_logic;
      dpc6: out std_logic;
      dpc7: out std_logic;
      dpc8: out std_logic;
      dpc9: out std_logic;
      dpc10: out std_logic;
      dpc11: out std_logic;
      dpc12: out std_logic;
      dpc13: out std_logic;
      ipc0: out std_logic;
      ipc1: out std_logic;
      ipc2: out std_logic;
      ipc3: out std_logic;
      ipc4: out std_logic;
      ipc5: out std_logic;
      ipc6: out std_logic;
      ipc7: out std_logic;
      ipc8: out std_logic;
      ipc9: out std_logic;
      ipc10: out std_logic;
      ipc11: out std_logic;
      ipc12: out std_logic;
      ipc13: out std_logic;
      pc0: out std_logic;
      pc1: out std_logic;
      pc2: out std_logic;
      pc3: out std_logic;
      pc4: out std_logic;
      pc5: out std_logic;
      pc6: out std_logic;
      pc7: out std_logic;
      pc8: out std_logic;
      pc9: out std_logic;
      pc10: out std_logic;
      pc11: out std_logic;
      pc12: out std_logic;
      pc13: out std_logic;
      spc0: out std_logic;
      spc2: out std_logic;
      spc3: out std_logic;
      spc4: out std_logic;
      spc5: out std_logic;
      spc6: out std_logic;
      spc7: out std_logic;
      spc8: out std_logic;
      spc9: out std_logic;
      spc10: out std_logic;
      spc11: out std_logic;
      spc12: out std_logic;
      spc13: out std_logic
    );
  end component;
  component olord_set is
      -- internal signals: \-boot\ \-clock reset a\ \-errhalt\ errstop mclk5a 
      -- internal signals: \stat.ovf\ statstop 
    port (
      aparok: in std_logic;
      clk5: in std_logic;
      dparok: in std_logic;
      iparok: in std_logic;
      \-ldclk\: in std_logic;
      \-ldopc\: in std_logic;
      mclk5: in std_logic;
      memparok: in std_logic;
      mmemparok: in std_logic;
      pdlparok: in std_logic;
      spcparok: in std_logic;
      spy0: in std_logic;
      spy1: in std_logic;
      spy2: in std_logic;
      spy3: in std_logic;
      spy4: in std_logic;
      spy5: in std_logic;
      spy6: in std_logic;
      spy7: in std_logic;
      \-stc32\: in std_logic;
      \-tpr60\: in std_logic;
      \-upperhighok\: in std_logic;
      v0parok: in std_logic;
      vmoparok: in std_logic;
      \-wait\: in std_logic;
      \-ldmode\: inout std_logic;
      \-reset\: inout std_logic;
      \-ape\: out std_logic;
      \boot.trap\: out std_logic;
      \-clk5\: out std_logic;
      clk5a: out std_logic;
      \-clock reset b\: out std_logic;
      \-dpe\: out std_logic;
      err: out std_logic;
      hi1: out std_logic;
      hi2: out std_logic;
      \-higherr\: out std_logic;
      idebug: out std_logic;
      \-idebug\: out std_logic;
      \-ipe\: out std_logic;
      \-ldstat\: out std_logic;
      \lpc.hold\: out std_logic;
      machrun: out std_logic;
      \-machruna\: out std_logic;
      \-mempe\: out std_logic;
      \-mpe\: out std_logic;
      \-nop11\: out std_logic;
      opcclk: out std_logic;
      \-opcinh\: out std_logic;
      \-pdlpe\: out std_logic;
      promdisable: out std_logic;
      promdisabled: out std_logic;
      reset: out std_logic;
      \-spe\: out std_logic;
      srun: out std_logic;
      ssdone: out std_logic;
      sspeed0: out std_logic;
      sspeed1: out std_logic;
      \-stathalt\: out std_logic;
      trapenb: out std_logic;
      \-v0pe\: out std_logic;
      \-v1pe\: out std_logic
    );
  end component;
  component opc_set is

    port (
      \-clk5\: in std_logic;
      dc0: in std_logic;
      dc1: in std_logic;
      dc2: in std_logic;
      dc3: in std_logic;
      dc4: in std_logic;
      dc5: in std_logic;
      dc6: in std_logic;
      dc7: in std_logic;
      dc8: in std_logic;
      dc9: in std_logic;
      hi2: in std_logic;
      opcclk: in std_logic;
      \-opcinh\: in std_logic;
      pc0: in std_logic;
      pc1: in std_logic;
      pc2: in std_logic;
      pc3: in std_logic;
      pc4: in std_logic;
      pc5: in std_logic;
      pc6: in std_logic;
      pc7: in std_logic;
      pc8: in std_logic;
      pc9: in std_logic;
      pc10: in std_logic;
      pc11: in std_logic;
      pc12: in std_logic;
      pc13: in std_logic;
      \-srcdc\: in std_logic;
      \-srcopc\: in std_logic;
      \-srcpdlidx\: in std_logic;
      \-srcpdlptr\: in std_logic;
      tse1b: in std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mf12: out std_logic;
      mf13: out std_logic;
      mf14: out std_logic;
      mf15: out std_logic;
      mf16: out std_logic;
      mf17: out std_logic;
      mf18: out std_logic;
      mf19: out std_logic;
      mf20: out std_logic;
      mf21: out std_logic;
      mf22: out std_logic;
      mf23: out std_logic;
      mf24: out std_logic;
      mf25: out std_logic;
      mf26: out std_logic;
      mf27: out std_logic;
      mf28: out std_logic;
      mf29: out std_logic;
      mf30: out std_logic;
      mf31: out std_logic;
      opc0: out std_logic;
      opc1: out std_logic;
      opc2: out std_logic;
      opc3: out std_logic;
      opc4: out std_logic;
      opc5: out std_logic;
      opc6: out std_logic;
      opc7: out std_logic;
      opc8: out std_logic;
      opc9: out std_logic;
      opc10: out std_logic;
      opc11: out std_logic;
      opc12: out std_logic;
      opc13: out std_logic
    );
  end component;
  component pdl_set is
      -- internal signals: pdl0 pdl1 pdl2 pdl3 pdl4 
      -- internal signals: pdl5 pdl6 pdl7 pdl8 pdl9 
      -- internal signals: pdl10 pdl11 pdl12 pdl13 pdl14 
      -- internal signals: pdl15 pdl16 pdl17 pdl18 pdl19 
      -- internal signals: pdl20 pdl21 pdl22 pdl23 pdl24 
      -- internal signals: pdl25 pdl26 pdl27 pdl28 pdl29 
      -- internal signals: pdl30 pdl31 \-pdla0a\ \-pdla0b\ \-pdla1a\ 
      -- internal signals: \-pdla1b\ \-pdla2a\ \-pdla2b\ \-pdla3a\ \-pdla3b\ 
      -- internal signals: \-pdla4a\ \-pdla4b\ \-pdla5a\ \-pdla5b\ \-pdla6a\ 
      -- internal signals: \-pdla6b\ \-pdla7a\ \-pdla7b\ \-pdla8a\ \-pdla8b\ 
      -- internal signals: \-pdla9a\ \-pdla9b\ \-pdlcnt\ \-pdldrive\ pdlidx0 
      -- internal signals: pdlidx1 pdlidx2 pdlidx3 pdlidx4 pdlidx5 
      -- internal signals: pdlidx6 pdlidx7 pdlidx8 pdlidx9 pdlparity 
      -- internal signals: pdlptr0 pdlptr1 pdlptr2 pdlptr3 pdlptr4 
      -- internal signals: pdlptr5 pdlptr6 pdlptr7 pdlptr8 pdlptr9 
      -- internal signals: \-pwpa\ \-pwpb\ \-pwpc\ 
    port (
      clk3f: in std_logic;
      clk4a: in std_logic;
      clk4b: in std_logic;
      clk4f: in std_logic;
      \-clk4e\: in std_logic;
      \-destpdl(p)\: in std_logic;
      \-destpdl(x)\: in std_logic;
      \-destpdlp\: in std_logic;
      \-destpdltop\: in std_logic;
      \-destpdlx\: in std_logic;
      \-destspc\: in std_logic;
      imod: in std_logic;
      ir30: in std_logic;
      l0: in std_logic;
      l1: in std_logic;
      l2: in std_logic;
      l3: in std_logic;
      l4: in std_logic;
      l5: in std_logic;
      l6: in std_logic;
      l7: in std_logic;
      l8: in std_logic;
      l9: in std_logic;
      l10: in std_logic;
      l11: in std_logic;
      l12: in std_logic;
      l13: in std_logic;
      l14: in std_logic;
      l15: in std_logic;
      l16: in std_logic;
      l17: in std_logic;
      l18: in std_logic;
      l19: in std_logic;
      l20: in std_logic;
      l21: in std_logic;
      l22: in std_logic;
      l23: in std_logic;
      l24: in std_logic;
      l25: in std_logic;
      l26: in std_logic;
      l27: in std_logic;
      l28: in std_logic;
      l29: in std_logic;
      l30: in std_logic;
      l31: in std_logic;
      lparity: in std_logic;
      nop: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      \-reset\: in std_logic;
      srcpdlidx: in std_logic;
      \-srcpdlpop\: in std_logic;
      srcpdlptr: in std_logic;
      \-srcpdltop\: in std_logic;
      tse4b: in std_logic;
      wp4a: in std_logic;
      imodd: out std_logic;
      m0: out std_logic;
      m1: out std_logic;
      m2: out std_logic;
      m3: out std_logic;
      m4: out std_logic;
      m5: out std_logic;
      m6: out std_logic;
      m7: out std_logic;
      m8: out std_logic;
      m9: out std_logic;
      m10: out std_logic;
      m11: out std_logic;
      m12: out std_logic;
      m13: out std_logic;
      m14: out std_logic;
      m15: out std_logic;
      m16: out std_logic;
      m17: out std_logic;
      m18: out std_logic;
      m19: out std_logic;
      m20: out std_logic;
      m21: out std_logic;
      m22: out std_logic;
      m23: out std_logic;
      m24: out std_logic;
      m25: out std_logic;
      m26: out std_logic;
      m27: out std_logic;
      m28: out std_logic;
      m29: out std_logic;
      m30: out std_logic;
      m31: out std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mparity: out std_logic;
      pdlenb: out std_logic;
      pdlwrited: out std_logic
    );
  end component;
  component prom_set is
      -- internal signals: \-promce0\ \-promce1\ \-prompc0\ \-prompc1\ \-prompc2\ 
      -- internal signals: \-prompc3\ \-prompc4\ \-prompc5\ \-prompc6\ \-prompc7\ 
      -- internal signals: \-prompc8\ 
    port (
      \-ape\: in std_logic;
      \-dpe\: in std_logic;
      hi2: in std_logic;
      \-idebug\: in std_logic;
      \-ipe\: in std_logic;
      \-iwriteda\: in std_logic;
      \-mempe\: in std_logic;
      \-mpe\: in std_logic;
      pc0: in std_logic;
      pc1: in std_logic;
      pc2: in std_logic;
      pc3: in std_logic;
      pc4: in std_logic;
      pc5: in std_logic;
      pc6: in std_logic;
      pc7: in std_logic;
      pc8: in std_logic;
      pc9: in std_logic;
      pc10: in std_logic;
      pc11: in std_logic;
      pc12: in std_logic;
      pc13: in std_logic;
      \-pdlpe\: in std_logic;
      \-promdisabled\: in std_logic;
      \-spe\: in std_logic;
      \-v0pe\: in std_logic;
      \-v1pe\: in std_logic;
      i0: out std_logic;
      i1: out std_logic;
      i2: out std_logic;
      i3: out std_logic;
      i4: out std_logic;
      i5: out std_logic;
      i6: out std_logic;
      i7: out std_logic;
      i8: out std_logic;
      i9: out std_logic;
      i10: out std_logic;
      i11: out std_logic;
      i12: out std_logic;
      i13: out std_logic;
      i14: out std_logic;
      i15: out std_logic;
      i16: out std_logic;
      i17: out std_logic;
      i18: out std_logic;
      i19: out std_logic;
      i20: out std_logic;
      i21: out std_logic;
      i22: out std_logic;
      i23: out std_logic;
      i24: out std_logic;
      i25: out std_logic;
      i26: out std_logic;
      i27: out std_logic;
      i28: out std_logic;
      i29: out std_logic;
      i30: out std_logic;
      i31: out std_logic;
      i32: out std_logic;
      i33: out std_logic;
      i34: out std_logic;
      i35: out std_logic;
      i36: out std_logic;
      i37: out std_logic;
      i38: out std_logic;
      i39: out std_logic;
      i40: out std_logic;
      i41: out std_logic;
      i42: out std_logic;
      i43: out std_logic;
      i44: out std_logic;
      i45: out std_logic;
      i46: out std_logic;
      i47: out std_logic;
      i48: out std_logic
    );
  end component;
  component qreg_set is
      -- internal signals: \-alu31\ q1 q2 q3 q4 
      -- internal signals: q5 q6 q7 q8 q9 
      -- internal signals: q10 q11 q12 q13 q14 
      -- internal signals: q15 q16 q17 q18 q19 
      -- internal signals: q20 q21 q22 q23 q24 
      -- internal signals: q25 q26 q27 q28 q29 
      -- internal signals: q30 qs0 qs1 
    port (
      alu0: in std_logic;
      alu1: in std_logic;
      alu2: in std_logic;
      alu3: in std_logic;
      alu4: in std_logic;
      alu5: in std_logic;
      alu6: in std_logic;
      alu7: in std_logic;
      alu8: in std_logic;
      alu9: in std_logic;
      alu10: in std_logic;
      alu11: in std_logic;
      alu12: in std_logic;
      alu13: in std_logic;
      alu14: in std_logic;
      alu15: in std_logic;
      alu16: in std_logic;
      alu17: in std_logic;
      alu18: in std_logic;
      alu19: in std_logic;
      alu20: in std_logic;
      alu21: in std_logic;
      alu22: in std_logic;
      alu23: in std_logic;
      alu24: in std_logic;
      alu25: in std_logic;
      alu26: in std_logic;
      alu27: in std_logic;
      alu28: in std_logic;
      alu29: in std_logic;
      alu30: in std_logic;
      alu31: in std_logic;
      clk2b: in std_logic;
      hi7: in std_logic;
      \-ir0\: in std_logic;
      \-ir1\: in std_logic;
      \-iralu\: in std_logic;
      \-srcq\: in std_logic;
      tse2: in std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mf12: out std_logic;
      mf13: out std_logic;
      mf14: out std_logic;
      mf15: out std_logic;
      mf16: out std_logic;
      mf17: out std_logic;
      mf18: out std_logic;
      mf19: out std_logic;
      mf20: out std_logic;
      mf21: out std_logic;
      mf22: out std_logic;
      mf23: out std_logic;
      mf24: out std_logic;
      mf25: out std_logic;
      mf26: out std_logic;
      mf27: out std_logic;
      mf28: out std_logic;
      mf29: out std_logic;
      mf30: out std_logic;
      mf31: out std_logic;
      q0: out std_logic;
      q31: out std_logic
    );
  end component;
  component shifter_masker_set is
      -- internal signals: mskl0 mskl1 mskl2 mskl3 mskl4 
      -- internal signals: mskr0 mskr1 mskr2 mskr3 mskr4 
      -- internal signals: s0 s1 s4 s2a s2b 
      -- internal signals: s3a s3b \-s4\ sa0 sa1 
      -- internal signals: sa2 sa3 sa4 sa5 sa6 
      -- internal signals: sa7 sa8 sa9 sa10 sa11 
      -- internal signals: sa12 sa13 sa14 sa15 sa16 
      -- internal signals: sa17 sa18 sa19 sa20 sa21 
      -- internal signals: sa22 sa23 sa24 sa25 sa26 
      -- internal signals: sa27 sa28 sa29 sa30 sa31 
    port (
      ir5: in std_logic;
      ir6: in std_logic;
      ir7: in std_logic;
      ir8: in std_logic;
      ir9: in std_logic;
      \-ir0\: in std_logic;
      ir12: in std_logic;
      ir13: in std_logic;
      \-ir1\: in std_logic;
      \-ir2\: in std_logic;
      ir31: in std_logic;
      \-irbyte\: in std_logic;
      m0: in std_logic;
      m1: in std_logic;
      m2: in std_logic;
      m3: in std_logic;
      m4: in std_logic;
      m6: in std_logic;
      m7: in std_logic;
      m8: in std_logic;
      m9: in std_logic;
      m10: in std_logic;
      m11: in std_logic;
      m12: in std_logic;
      m13: in std_logic;
      m14: in std_logic;
      m15: in std_logic;
      m16: in std_logic;
      m17: in std_logic;
      m18: in std_logic;
      m19: in std_logic;
      m20: in std_logic;
      m21: in std_logic;
      m22: in std_logic;
      m23: in std_logic;
      m24: in std_logic;
      m25: in std_logic;
      m26: in std_logic;
      m27: in std_logic;
      m28: in std_logic;
      m29: in std_logic;
      m30: in std_logic;
      m31: in std_logic;
      \-sh3\: in std_logic;
      \-sh4\: in std_logic;
      \a=m\: out std_logic;
      \-ir12\: out std_logic;
      \-ir13\: out std_logic;
      \-ir31\: out std_logic;
      m5: out std_logic;
      msk0: out std_logic;
      msk1: out std_logic;
      msk2: out std_logic;
      msk3: out std_logic;
      msk4: out std_logic;
      msk5: out std_logic;
      msk6: out std_logic;
      msk7: out std_logic;
      msk8: out std_logic;
      msk9: out std_logic;
      msk10: out std_logic;
      msk11: out std_logic;
      msk12: out std_logic;
      msk13: out std_logic;
      msk14: out std_logic;
      msk15: out std_logic;
      msk16: out std_logic;
      msk17: out std_logic;
      msk18: out std_logic;
      msk19: out std_logic;
      msk20: out std_logic;
      msk21: out std_logic;
      msk22: out std_logic;
      msk23: out std_logic;
      msk24: out std_logic;
      msk25: out std_logic;
      msk26: out std_logic;
      msk27: out std_logic;
      msk28: out std_logic;
      msk29: out std_logic;
      msk30: out std_logic;
      msk31: out std_logic;
      r0: out std_logic;
      r1: out std_logic;
      r2: out std_logic;
      r3: out std_logic;
      r4: out std_logic;
      r5: out std_logic;
      r6: out std_logic;
      r7: out std_logic;
      r8: out std_logic;
      r9: out std_logic;
      r10: out std_logic;
      r11: out std_logic;
      r12: out std_logic;
      r13: out std_logic;
      r14: out std_logic;
      r15: out std_logic;
      r16: out std_logic;
      r17: out std_logic;
      r18: out std_logic;
      r19: out std_logic;
      r20: out std_logic;
      r21: out std_logic;
      r22: out std_logic;
      r23: out std_logic;
      r24: out std_logic;
      r25: out std_logic;
      r26: out std_logic;
      r27: out std_logic;
      r28: out std_logic;
      r29: out std_logic;
      r30: out std_logic;
      r31: out std_logic
    );
  end component;
  component spc_set is
      -- internal signals: spc15 spc16 spc17 spc18 spco0 
      -- internal signals: spco1 spco2 spco3 spco4 spco5 
      -- internal signals: spco6 spco7 spco8 spco9 spco10 
      -- internal signals: spco11 spco12 spco13 spco14 spco15 
      -- internal signals: spco16 spco17 spco18 spcopar spcpar 
      -- internal signals: spcptr0 spcptr1 spcptr2 spcptr3 spcptr4 
      -- internal signals: spcw0 spcw1 spcw2 spcw3 spcw4 
      -- internal signals: spcw5 spcw6 spcw7 spcw8 spcw9 
      -- internal signals: spcw10 spcw11 spcw12 spcw13 spcw14 
      -- internal signals: spcw15 spcw16 spcw17 spcw18 spcwpar 
      -- internal signals: wpc0 wpc1 wpc2 wpc3 wpc4 
      -- internal signals: wpc5 wpc6 wpc7 wpc8 wpc9 
      -- internal signals: wpc10 wpc11 wpc12 wpc13 
    port (
      clk4b: in std_logic;
      clk4c: in std_logic;
      clk4d: in std_logic;
      clk4f: in std_logic;
      destspcd: in std_logic;
      ipc0: in std_logic;
      ipc1: in std_logic;
      ipc2: in std_logic;
      ipc3: in std_logic;
      ipc4: in std_logic;
      ipc5: in std_logic;
      ipc6: in std_logic;
      ipc7: in std_logic;
      ipc8: in std_logic;
      ipc9: in std_logic;
      ipc10: in std_logic;
      ipc11: in std_logic;
      ipc12: in std_logic;
      ipc13: in std_logic;
      ir25: in std_logic;
      irdisp: in std_logic;
      l0: in std_logic;
      l1: in std_logic;
      l2: in std_logic;
      l3: in std_logic;
      l4: in std_logic;
      l5: in std_logic;
      l6: in std_logic;
      l7: in std_logic;
      l8: in std_logic;
      l9: in std_logic;
      l10: in std_logic;
      l11: in std_logic;
      l12: in std_logic;
      l13: in std_logic;
      l14: in std_logic;
      l15: in std_logic;
      l16: in std_logic;
      l17: in std_logic;
      l18: in std_logic;
      \lpc.hold\: in std_logic;
      n: in std_logic;
      pc0: in std_logic;
      pc1: in std_logic;
      pc2: in std_logic;
      pc3: in std_logic;
      pc4: in std_logic;
      pc5: in std_logic;
      pc6: in std_logic;
      pc7: in std_logic;
      pc8: in std_logic;
      pc9: in std_logic;
      pc10: in std_logic;
      pc11: in std_logic;
      pc12: in std_logic;
      pc13: in std_logic;
      spcdrive: in std_logic;
      \-spcdrive\: in std_logic;
      \-spcnt\: in std_logic;
      \-spcpass\: in std_logic;
      spcwpass: in std_logic;
      \-spcwpass\: in std_logic;
      spush: in std_logic;
      \-swpa\: in std_logic;
      \-swpb\: in std_logic;
      hi1: inout std_logic;
      spc0: inout std_logic;
      spc2: inout std_logic;
      spc3: inout std_logic;
      spc4: inout std_logic;
      spc5: inout std_logic;
      spc6: inout std_logic;
      spc7: inout std_logic;
      spc8: inout std_logic;
      spc9: inout std_logic;
      spc10: inout std_logic;
      spc11: inout std_logic;
      spc12: inout std_logic;
      spc13: inout std_logic;
      hi2: out std_logic;
      hi3: out std_logic;
      hi4: out std_logic;
      hi5: out std_logic;
      hi6: out std_logic;
      hi7: out std_logic;
      hi8: out std_logic;
      hi9: out std_logic;
      hi10: out std_logic;
      hi11: out std_logic;
      hi12: out std_logic;
      m0: out std_logic;
      m1: out std_logic;
      m2: out std_logic;
      m3: out std_logic;
      m4: out std_logic;
      m5: out std_logic;
      m6: out std_logic;
      m7: out std_logic;
      m8: out std_logic;
      m9: out std_logic;
      m10: out std_logic;
      m11: out std_logic;
      m12: out std_logic;
      m13: out std_logic;
      m14: out std_logic;
      m15: out std_logic;
      m16: out std_logic;
      m17: out std_logic;
      m18: out std_logic;
      m19: out std_logic;
      m20: out std_logic;
      m21: out std_logic;
      m22: out std_logic;
      m23: out std_logic;
      m24: out std_logic;
      m25: out std_logic;
      m26: out std_logic;
      m27: out std_logic;
      m28: out std_logic;
      m29: out std_logic;
      m30: out std_logic;
      m31: out std_logic;
      spc1: out std_logic;
      spc14: out std_logic;
      spcparok: out std_logic
    );
  end component;
  component spy_set is
      -- internal signals: \-spy.ah\ \-spy.flag2\ \-spy.irh\ \-spy.irl\ \-spy.irm\ 
      -- internal signals: \-spy.mh\ \-spy.ml\ \-spy.obh\ \-spy.opc\ \-spy.pc\ 
    port (
      a16: in std_logic;
      a17: in std_logic;
      a18: in std_logic;
      a19: in std_logic;
      a20: in std_logic;
      a21: in std_logic;
      a22: in std_logic;
      a23: in std_logic;
      a24: in std_logic;
      a25: in std_logic;
      a26: in std_logic;
      a27: in std_logic;
      a28: in std_logic;
      a29: in std_logic;
      a30: in std_logic;
      a31a: in std_logic;
      aa0: in std_logic;
      aa1: in std_logic;
      aa2: in std_logic;
      aa3: in std_logic;
      aa4: in std_logic;
      aa5: in std_logic;
      aa6: in std_logic;
      aa7: in std_logic;
      aa8: in std_logic;
      aa9: in std_logic;
      aa10: in std_logic;
      aa11: in std_logic;
      aa12: in std_logic;
      aa13: in std_logic;
      aa14: in std_logic;
      aa15: in std_logic;
      \-ape\: in std_logic;
      destspcd: in std_logic;
      \-dpe\: in std_logic;
      err: in std_logic;
      hi1: in std_logic;
      \-higherr\: in std_logic;
      imodd: in std_logic;
      \-ipe\: in std_logic;
      ir0: in std_logic;
      ir1: in std_logic;
      ir2: in std_logic;
      ir3: in std_logic;
      ir4: in std_logic;
      ir5: in std_logic;
      ir6: in std_logic;
      ir7: in std_logic;
      ir8: in std_logic;
      ir9: in std_logic;
      ir10: in std_logic;
      ir11: in std_logic;
      ir12: in std_logic;
      ir13: in std_logic;
      ir14: in std_logic;
      ir15: in std_logic;
      ir16: in std_logic;
      ir17: in std_logic;
      ir18: in std_logic;
      ir19: in std_logic;
      ir20: in std_logic;
      ir21: in std_logic;
      ir22: in std_logic;
      ir23: in std_logic;
      ir24: in std_logic;
      ir25: in std_logic;
      ir26: in std_logic;
      ir27: in std_logic;
      ir28: in std_logic;
      ir29: in std_logic;
      ir30: in std_logic;
      ir31: in std_logic;
      ir32: in std_logic;
      ir33: in std_logic;
      ir34: in std_logic;
      ir35: in std_logic;
      ir36: in std_logic;
      ir37: in std_logic;
      ir38: in std_logic;
      ir39: in std_logic;
      ir40: in std_logic;
      ir41: in std_logic;
      ir42: in std_logic;
      ir43: in std_logic;
      ir44: in std_logic;
      ir45: in std_logic;
      ir46: in std_logic;
      ir47: in std_logic;
      ir48: in std_logic;
      iwrited: in std_logic;
      jcond: in std_logic;
      m0: in std_logic;
      m1: in std_logic;
      m2: in std_logic;
      m3: in std_logic;
      m4: in std_logic;
      m5: in std_logic;
      m6: in std_logic;
      m7: in std_logic;
      m8: in std_logic;
      m9: in std_logic;
      m10: in std_logic;
      m11: in std_logic;
      m12: in std_logic;
      m13: in std_logic;
      m14: in std_logic;
      m15: in std_logic;
      m16: in std_logic;
      m17: in std_logic;
      m18: in std_logic;
      m19: in std_logic;
      m20: in std_logic;
      m21: in std_logic;
      m22: in std_logic;
      m23: in std_logic;
      m24: in std_logic;
      m25: in std_logic;
      m26: in std_logic;
      m27: in std_logic;
      m28: in std_logic;
      m29: in std_logic;
      m30: in std_logic;
      m31: in std_logic;
      \-mempe\: in std_logic;
      \-mpe\: in std_logic;
      nop: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      ob10: in std_logic;
      ob11: in std_logic;
      ob12: in std_logic;
      ob13: in std_logic;
      ob14: in std_logic;
      ob15: in std_logic;
      ob16: in std_logic;
      ob17: in std_logic;
      ob18: in std_logic;
      ob19: in std_logic;
      ob20: in std_logic;
      ob21: in std_logic;
      ob22: in std_logic;
      ob23: in std_logic;
      ob24: in std_logic;
      ob25: in std_logic;
      ob26: in std_logic;
      ob27: in std_logic;
      ob28: in std_logic;
      ob29: in std_logic;
      ob30: in std_logic;
      ob31: in std_logic;
      opc0: in std_logic;
      opc1: in std_logic;
      opc2: in std_logic;
      opc3: in std_logic;
      opc4: in std_logic;
      opc5: in std_logic;
      opc6: in std_logic;
      opc7: in std_logic;
      opc8: in std_logic;
      opc9: in std_logic;
      opc10: in std_logic;
      opc11: in std_logic;
      opc12: in std_logic;
      opc13: in std_logic;
      pc0: in std_logic;
      pc1: in std_logic;
      pc2: in std_logic;
      pc3: in std_logic;
      pc4: in std_logic;
      pc5: in std_logic;
      pc6: in std_logic;
      pc7: in std_logic;
      pc8: in std_logic;
      pc9: in std_logic;
      pc10: in std_logic;
      pc11: in std_logic;
      pc12: in std_logic;
      pc13: in std_logic;
      pcs0: in std_logic;
      pcs1: in std_logic;
      \-pdlpe\: in std_logic;
      pdlwrited: in std_logic;
      promdisable: in std_logic;
      \-spe\: in std_logic;
      spushd: in std_logic;
      srun: in std_logic;
      ssdone: in std_logic;
      \-stathalt\: in std_logic;
      \-v0pe\: in std_logic;
      \-v1pe\: in std_logic;
      \-vmaok\: in std_logic;
      \-wait\: in std_logic;
      wmapd: in std_logic;
      \-ldclk\: out std_logic;
      \-lddbirh\: out std_logic;
      \-lddbirl\: out std_logic;
      \-lddbirm\: out std_logic;
      \-ldmode\: out std_logic;
      \-ldopc\: out std_logic;
      \-spy.sth\: out std_logic;
      \-spy.stl\: out std_logic;
      spy0: out std_logic;
      spy1: out std_logic;
      spy2: out std_logic;
      spy3: out std_logic;
      spy4: out std_logic;
      spy5: out std_logic;
      spy6: out std_logic;
      spy7: out std_logic;
      spy8: out std_logic;
      spy9: out std_logic;
      spy10: out std_logic;
      spy11: out std_logic;
      spy12: out std_logic;
      spy13: out std_logic;
      spy14: out std_logic;
      spy15: out std_logic
    );
  end component;
  component stat_set is

    port (
      clk5a: in std_logic;
      hi1: in std_logic;
      iwr0: in std_logic;
      iwr1: in std_logic;
      iwr2: in std_logic;
      iwr3: in std_logic;
      iwr4: in std_logic;
      iwr5: in std_logic;
      iwr6: in std_logic;
      iwr7: in std_logic;
      iwr8: in std_logic;
      iwr9: in std_logic;
      iwr10: in std_logic;
      iwr11: in std_logic;
      iwr12: in std_logic;
      iwr13: in std_logic;
      iwr14: in std_logic;
      iwr15: in std_logic;
      iwr16: in std_logic;
      iwr17: in std_logic;
      iwr18: in std_logic;
      iwr19: in std_logic;
      iwr20: in std_logic;
      iwr21: in std_logic;
      iwr22: in std_logic;
      iwr23: in std_logic;
      iwr24: in std_logic;
      iwr25: in std_logic;
      iwr26: in std_logic;
      iwr27: in std_logic;
      iwr28: in std_logic;
      iwr29: in std_logic;
      iwr30: in std_logic;
      iwr31: in std_logic;
      \-ldstat\: in std_logic;
      \-spy.sth\: in std_logic;
      \-spy.stl\: in std_logic;
      \-statbit\: in std_logic;
      spy0: out std_logic;
      spy1: out std_logic;
      spy2: out std_logic;
      spy3: out std_logic;
      spy4: out std_logic;
      spy5: out std_logic;
      spy6: out std_logic;
      spy7: out std_logic;
      spy8: out std_logic;
      spy9: out std_logic;
      spy10: out std_logic;
      spy11: out std_logic;
      spy12: out std_logic;
      spy13: out std_logic;
      spy14: out std_logic;
      spy15: out std_logic;
      \-stc32\: out std_logic
    );
  end component;
  component trap_set is

    port (
      \boot.trap\: in std_logic;
      \-md0\: in std_logic;
      \-md1\: in std_logic;
      \-md2\: in std_logic;
      \-md3\: in std_logic;
      \-md4\: in std_logic;
      \-md5\: in std_logic;
      \-md6\: in std_logic;
      \-md7\: in std_logic;
      \-md8\: in std_logic;
      \-md9\: in std_logic;
      \-md10\: in std_logic;
      \-md11\: in std_logic;
      \-md12\: in std_logic;
      \-md13\: in std_logic;
      \-md14\: in std_logic;
      \-md15\: in std_logic;
      \-md16\: in std_logic;
      \-md17\: in std_logic;
      \-md18\: in std_logic;
      \-md19\: in std_logic;
      \-md20\: in std_logic;
      \-md21\: in std_logic;
      \-md22\: in std_logic;
      \-md23\: in std_logic;
      \-md24\: in std_logic;
      \-md25\: in std_logic;
      \-md26\: in std_logic;
      \-md27\: in std_logic;
      \-md28\: in std_logic;
      \-md29\: in std_logic;
      \-md30\: in std_logic;
      \-md31\: in std_logic;
      mdhaspar: in std_logic;
      mdpar: in std_logic;
      trapenb: in std_logic;
      \use.md\: in std_logic;
      \-wait\: in std_logic;
      mdparodd: out std_logic;
      memparok: out std_logic;
      \-trap\: out std_logic;
      trapa: out std_logic;
      trapb: out std_logic
    );
  end component;
  component vctl_set is
      -- internal signals: destmem memprepare \-memprepare\ \-memrd\ memrq 
      -- internal signals: \-memwr\ wmap wrcyc 
    port (
      clk2a: in std_logic;
      clk2c: in std_logic;
      \-clk3g\: in std_logic;
      \-destmdr\: in std_logic;
      \-destmem\: in std_logic;
      \-destvma\: in std_logic;
      hi4: in std_logic;
      hi11: in std_logic;
      \-ifetch\: in std_logic;
      ir19: in std_logic;
      ir20: in std_logic;
      lcinc: in std_logic;
      \-lvmo22\: in std_logic;
      \-lvmo23\: in std_logic;
      mclk1a: in std_logic;
      needfetch: in std_logic;
      \-nopa\: in std_logic;
      \-reset\: in std_logic;
      \-srcmd\: in std_logic;
      \-vma25\: in std_logic;
      \-vma26\: in std_logic;
      wp1a: in std_logic;
      wp1b: in std_logic;
      \-hang\: out std_logic;
      mdsela: out std_logic;
      mdselb: out std_logic;
      \-memdrive.a\: out std_logic;
      \-memdrive.b\: out std_logic;
      memstart: out std_logic;
      \-memstart\: out std_logic;
      \-pfr\: out std_logic;
      \-pfw\: out std_logic;
      \use.md\: out std_logic;
      \-vm0wpa\: out std_logic;
      \-vm0wpb\: out std_logic;
      \-vm1wpa\: out std_logic;
      \-vm1wpb\: out std_logic;
      \-vmaenb\: out std_logic;
      \-vmaok\: out std_logic;
      vmasela: out std_logic;
      vmaselb: out std_logic;
      \-wait\: out std_logic;
      wmapd: out std_logic
    );
  end component;
  component vma_set is
      -- internal signals: \-vmas0\ \-vmas1\ \-vmas2\ \-vmas3\ \-vmas4\ 
      -- internal signals: \-vmas5\ \-vmas6\ \-vmas7\ \-vmas8\ \-vmas9\ 
      -- internal signals: \-vmas10\ \-vmas11\ \-vmas12\ \-vmas13\ \-vmas14\ 
      -- internal signals: \-vmas15\ \-vmas16\ \-vmas17\ \-vmas18\ \-vmas19\ 
      -- internal signals: \-vmas20\ \-vmas21\ \-vmas22\ \-vmas23\ \-vmas24\ 
      -- internal signals: \-vmas25\ \-vmas26\ \-vmas27\ \-vmas28\ \-vmas29\ 
      -- internal signals: \-vmas30\ \-vmas31\ 
    port (
      clk1a: in std_logic;
      clk2a: in std_logic;
      clk2c: in std_logic;
      lc2: in std_logic;
      lc3: in std_logic;
      lc4: in std_logic;
      lc5: in std_logic;
      lc6: in std_logic;
      lc7: in std_logic;
      lc8: in std_logic;
      lc9: in std_logic;
      lc10: in std_logic;
      lc11: in std_logic;
      lc12: in std_logic;
      lc13: in std_logic;
      lc14: in std_logic;
      lc15: in std_logic;
      lc16: in std_logic;
      lc17: in std_logic;
      lc18: in std_logic;
      lc19: in std_logic;
      lc20: in std_logic;
      lc21: in std_logic;
      lc22: in std_logic;
      lc23: in std_logic;
      lc24: in std_logic;
      lc25: in std_logic;
      \-md8\: in std_logic;
      \-md9\: in std_logic;
      \-md10\: in std_logic;
      \-md11\: in std_logic;
      \-md12\: in std_logic;
      \-md13\: in std_logic;
      \-md14\: in std_logic;
      \-md15\: in std_logic;
      \-md16\: in std_logic;
      \-md17\: in std_logic;
      \-md18\: in std_logic;
      \-md19\: in std_logic;
      \-md20\: in std_logic;
      \-md21\: in std_logic;
      \-md22\: in std_logic;
      \-md23\: in std_logic;
      \-memstart\: in std_logic;
      ob0: in std_logic;
      ob1: in std_logic;
      ob2: in std_logic;
      ob3: in std_logic;
      ob4: in std_logic;
      ob5: in std_logic;
      ob6: in std_logic;
      ob7: in std_logic;
      ob8: in std_logic;
      ob9: in std_logic;
      ob10: in std_logic;
      ob11: in std_logic;
      ob12: in std_logic;
      ob13: in std_logic;
      ob14: in std_logic;
      ob15: in std_logic;
      ob16: in std_logic;
      ob17: in std_logic;
      ob18: in std_logic;
      ob19: in std_logic;
      ob20: in std_logic;
      ob21: in std_logic;
      ob22: in std_logic;
      ob23: in std_logic;
      ob24: in std_logic;
      ob25: in std_logic;
      ob26: in std_logic;
      ob27: in std_logic;
      ob28: in std_logic;
      ob29: in std_logic;
      ob30: in std_logic;
      ob31: in std_logic;
      \-srcvma\: in std_logic;
      tse2: in std_logic;
      \-vmaenb\: in std_logic;
      vmasela: in std_logic;
      vmaselb: in std_logic;
      mapi8: out std_logic;
      mapi9: out std_logic;
      mapi10: out std_logic;
      mapi11: out std_logic;
      mapi12: out std_logic;
      mapi13: out std_logic;
      mapi14: out std_logic;
      mapi15: out std_logic;
      mapi16: out std_logic;
      mapi17: out std_logic;
      mapi18: out std_logic;
      mapi19: out std_logic;
      mapi20: out std_logic;
      mapi21: out std_logic;
      mapi22: out std_logic;
      mapi23: out std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mf12: out std_logic;
      mf13: out std_logic;
      mf14: out std_logic;
      mf15: out std_logic;
      mf16: out std_logic;
      mf17: out std_logic;
      mf18: out std_logic;
      mf19: out std_logic;
      mf20: out std_logic;
      mf21: out std_logic;
      mf22: out std_logic;
      mf23: out std_logic;
      mf24: out std_logic;
      mf25: out std_logic;
      mf26: out std_logic;
      mf27: out std_logic;
      mf28: out std_logic;
      mf29: out std_logic;
      mf30: out std_logic;
      mf31: out std_logic;
      \-vma0\: out std_logic;
      \-vma1\: out std_logic;
      \-vma2\: out std_logic;
      \-vma3\: out std_logic;
      \-vma4\: out std_logic;
      \-vma5\: out std_logic;
      \-vma6\: out std_logic;
      \-vma7\: out std_logic;
      \-vma8\: out std_logic;
      \-vma9\: out std_logic;
      \-vma10\: out std_logic;
      \-vma11\: out std_logic;
      \-vma12\: out std_logic;
      \-vma13\: out std_logic;
      \-vma14\: out std_logic;
      \-vma15\: out std_logic;
      \-vma16\: out std_logic;
      \-vma17\: out std_logic;
      \-vma18\: out std_logic;
      \-vma19\: out std_logic;
      \-vma20\: out std_logic;
      \-vma21\: out std_logic;
      \-vma22\: out std_logic;
      \-vma23\: out std_logic;
      \-vma25\: out std_logic;
      \-vma26\: out std_logic;
      \-vma27\: out std_logic;
      \-vma28\: out std_logic;
      \-vma29\: out std_logic;
      \-vma30\: out std_logic;
      \-vma31\: out std_logic
    );
  end component;
  component vmaps_set is
      -- internal signals: \-mapi8b\ \-mapi9b\ \-mapi10b\ \-mapi11b\ \-mapi12b\ 
      -- internal signals: srcmap vm1pari \-vmap0\ \-vmap1\ \-vmap2\ 
      -- internal signals: \-vmap3\ \-vmap4\ \-vmo0\ \-vmo1\ \-vmo2\ 
      -- internal signals: \-vmo3\ \-vmo4\ \-vmo5\ \-vmo6\ \-vmo7\ 
      -- internal signals: \-vmo8\ \-vmo9\ \-vmo10\ \-vmo11\ \-vmo12\ 
      -- internal signals: \-vmo13\ \-vmo14\ \-vmo15\ \-vmo16\ \-vmo17\ 
      -- internal signals: \-vmo20\ \-vmo21\ \-vmo22\ \-vmo23\ vmoparodd 
    port (
      hi12: in std_logic;
      mapi8: in std_logic;
      mapi9: in std_logic;
      mapi10: in std_logic;
      mapi11: in std_logic;
      mapi12: in std_logic;
      mapi13: in std_logic;
      mapi14: in std_logic;
      mapi15: in std_logic;
      mapi16: in std_logic;
      mapi17: in std_logic;
      mapi18: in std_logic;
      mapi19: in std_logic;
      mapi20: in std_logic;
      mapi21: in std_logic;
      mapi22: in std_logic;
      mapi23: in std_logic;
      memstart: in std_logic;
      \-pfr\: in std_logic;
      \-pfw\: in std_logic;
      \-srcmap\: in std_logic;
      tse1a: in std_logic;
      \-vm0wpa\: in std_logic;
      \-vm0wpb\: in std_logic;
      \-vm1wpa\: in std_logic;
      \-vm1wpb\: in std_logic;
      \-vma0\: in std_logic;
      \-vma1\: in std_logic;
      \-vma2\: in std_logic;
      \-vma3\: in std_logic;
      \-vma4\: in std_logic;
      \-vma5\: in std_logic;
      \-vma6\: in std_logic;
      \-vma7\: in std_logic;
      \-vma8\: in std_logic;
      \-vma9\: in std_logic;
      \-vma10\: in std_logic;
      \-vma11\: in std_logic;
      \-vma12\: in std_logic;
      \-vma13\: in std_logic;
      \-vma14\: in std_logic;
      \-vma15\: in std_logic;
      \-vma16\: in std_logic;
      \-vma17\: in std_logic;
      \-vma18\: in std_logic;
      \-vma19\: in std_logic;
      \-vma20\: in std_logic;
      \-vma21\: in std_logic;
      \-vma22\: in std_logic;
      \-vma23\: in std_logic;
      \-vma27\: in std_logic;
      \-vma28\: in std_logic;
      \-vma29\: in std_logic;
      \-vma30\: in std_logic;
      \-vma31\: in std_logic;
      \-vmo18\: inout std_logic;
      \-vmo19\: inout std_logic;
      \-lvmo22\: out std_logic;
      \-lvmo23\: out std_logic;
      mf0: out std_logic;
      mf1: out std_logic;
      mf2: out std_logic;
      mf3: out std_logic;
      mf4: out std_logic;
      mf5: out std_logic;
      mf6: out std_logic;
      mf7: out std_logic;
      mf8: out std_logic;
      mf9: out std_logic;
      mf10: out std_logic;
      mf11: out std_logic;
      mf12: out std_logic;
      mf13: out std_logic;
      mf14: out std_logic;
      mf15: out std_logic;
      mf16: out std_logic;
      mf17: out std_logic;
      mf18: out std_logic;
      mf19: out std_logic;
      mf20: out std_logic;
      mf21: out std_logic;
      mf22: out std_logic;
      mf23: out std_logic;
      mf24: out std_logic;
      mf25: out std_logic;
      mf26: out std_logic;
      mf27: out std_logic;
      mf28: out std_logic;
      mf29: out std_logic;
      mf30: out std_logic;
      mf31: out std_logic;
      v0parok: out std_logic;
      vmoparok: out std_logic
    );
  end component;
end package;
