library ieee;
use ieee.std_logic_1164.all;

entity cadr_vmem2 is
  port (
    \-mapi10b\      : in     std_logic;
    \-mapi11b\      : in     std_logic;
    \-mapi12b\      : in     std_logic;
    \-mapi8b\       : in     std_logic;
    \-mapi9b\       : in     std_logic;
    \-vm1wpb\       : in     std_logic;
    \-vma12\        : in     std_logic;
    \-vma13\        : in     std_logic;
    \-vma14\        : in     std_logic;
    \-vma15\        : in     std_logic;
    \-vma16\        : in     std_logic;
    \-vma17\        : in     std_logic;
    \-vma18\        : in     std_logic;
    \-vma19\        : in     std_logic;
    \-vma20\        : in     std_logic;
    \-vma21\        : in     std_logic;
    \-vma22\        : in     std_logic;
    \-vma23\        : in     std_logic;
    \-vmap0\        : in     std_logic;
    \-vmap1\        : in     std_logic;
    \-vmap2\        : in     std_logic;
    \-vmap3\        : in     std_logic;
    \-vmap4\        : in     std_logic;
    \-vmo0\         : in     std_logic;
    \-vmo10\        : in     std_logic;
    \-vmo11\        : in     std_logic;
    \-vmo1\         : in     std_logic;
    \-vmo2\         : in     std_logic;
    \-vmo3\         : in     std_logic;
    \-vmo4\         : in     std_logic;
    \-vmo5\         : in     std_logic;
    \-vmo6\         : in     std_logic;
    \-vmo7\         : in     std_logic;
    \-vmo8\         : in     std_logic;
    \-vmo9\         : in     std_logic;
    vm1pari         : in     std_logic;
    \-vmo12\        : out    std_logic;
    \-vmo13\        : out    std_logic;
    \-vmo14\        : out    std_logic;
    \-vmo15\        : out    std_logic;
    \-vmo16\        : out    std_logic;
    \-vmo17\        : out    std_logic;
    \-vmo18\        : out    std_logic;
    \-vmo19\        : out    std_logic;
    \-vmo20\        : out    std_logic;
    \-vmo21\        : out    std_logic;
    \-vmo22\        : out    std_logic;
    \-vmo23\        : out    std_logic;
    vmap0b          : out    std_logic;
    vmap1b          : out    std_logic;
    vmap2b          : out    std_logic;
    vmap3b          : out    std_logic;
    vmap4b          : out    std_logic;
    vmopar          : out    std_logic;
    vmoparck        : out    std_logic;
    vmoparl         : out    std_logic;
    vmoparm         : out    std_logic;
    vmoparodd       : out    std_logic
  );
end entity;
