-- 4 Bit Binary Full Adders With Fast Carry

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sn74283 is
  port (
    ci : in std_logic := 'H'; -- Pin 7
    a0 : in std_logic := 'H'; -- Pin 5
    a1 : in std_logic := 'H'; -- Pin 3
    a2 : in std_logic := 'H'; -- Pin 14
    a3 : in std_logic := 'H'; -- Pin 13
    b0 : in std_logic := 'H'; -- Pin 6
    b1 : in std_logic := 'H'; -- Pin 2
    b2 : in std_logic := 'H'; -- Pin 15
    b3 : in std_logic := 'H'; -- Pin 11
    s0 : out std_logic; -- Pin 4
    s1 : out std_logic; -- Pin 1
    s2 : out std_logic; -- Pin 13
    s3 : out std_logic; -- Pin 10
    co : out std_logic  -- Pin 9
    );
end;

architecture ttl of sn74283 is
  signal a : unsigned(3 downto 0);
  signal b : unsigned(3 downto 0);
begin
  a <= a3 & a2 & a1 & a0;
  b <= b3 & b2 & b1 & b0;

  process(all)
    variable sum : unsigned(4 downto 0);
  begin
    -- Check for unknown inputs
    if is_x(a) or is_x(b) then
      -- Any unknown input causes unknown outputs
      s0 <= 'X'; s1 <= 'X'; s2 <= 'X'; s3 <= 'X'; co <= 'X';
    else
      -- All inputs are valid, perform addition
      sum := ('0' & a) + ('0' & b) + ("0000" & ci);
      s3  <= sum(3); s2 <= sum(2); s1 <= sum(1); s0 <= sum(0);
      co  <= sum(4);
    end if;
  end process;
end;
