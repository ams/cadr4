library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_res20 is
  port (
    r2  : out std_logic;
    r3  : out std_logic;
    r4  : out std_logic;
    r5  : out std_logic;
    r6  : out std_logic;
    r7  : out std_logic;
    r8  : out std_logic;
    r9  : out std_logic;
    r10 : out std_logic;
    r11 : out std_logic;
    r12 : out std_logic;
    r13 : out std_logic;
    r14 : out std_logic;
    r15 : out std_logic;
    r16 : out std_logic;
    r17 : out std_logic;
    r18 : out std_logic;
    r19 : out std_logic
    );
end ic_res20;

architecture ttl of ic_res20 is
begin

end ttl;
