-- CADR1_UBMAP
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_ubmap is
  port (
    \-ubmap _ udo\ : in std_logic;
    \-ubmapwe\ : inout std_logic;
    \-ubpn0a\ : inout std_logic;
    \-ubpn0b\ : out std_logic;
    \-ubpn1a\ : inout std_logic;
    \-ubpn1b\ : out std_logic;
    \-ubpn2a\ : inout std_logic;
    \-ubpn2b\ : out std_logic;
    \-ubpn3a\ : inout std_logic;
    \-ubpn3b\ : out std_logic;
    mapvalid : inout std_logic;
    \select page\ : in std_logic;
    uba1 : in std_logic;
    uba10 : in std_logic;
    uba11 : in std_logic;
    uba12 : in std_logic;
    uba13 : in std_logic;
    uba2 : in std_logic;
    uba3 : in std_logic;
    uba4 : in std_logic;
    \ubma 10\ : in std_logic;
    \ubma 11\ : in std_logic;
    \ubma 12\ : in std_logic;
    \ubma 13\ : in std_logic;
    \ubma 14\ : in std_logic;
    \ubma 15\ : in std_logic;
    \ubma 16\ : in std_logic;
    \ubma 17\ : in std_logic;
    \ubma 18\ : in std_logic;
    \ubma 19\ : in std_logic;
    \ubma 20\ : in std_logic;
    \ubma 21\ : in std_logic;
    \ubma 8\ : in std_logic;
    \ubma 9\ : in std_logic;
    ubma10 : inout std_logic;
    ubma11 : inout std_logic;
    ubma12 : inout std_logic;
    ubma13 : inout std_logic;
    ubma14 : inout std_logic;
    ubma15 : inout std_logic;
    ubma16 : inout std_logic;
    ubma17 : inout std_logic;
    ubma18 : inout std_logic;
    ubma19 : inout std_logic;
    ubma20 : inout std_logic;
    ubma21 : inout std_logic;
    ubma8 : inout std_logic;
    ubma9 : inout std_logic;
    udi0 : inout std_logic;
    udi1 : inout std_logic;
    udi10 : inout std_logic;
    udi11 : inout std_logic;
    udi12 : inout std_logic;
    udi13 : inout std_logic;
    udi14 : inout std_logic;
    udi15 : inout std_logic;
    udi2 : inout std_logic;
    udi3 : inout std_logic;
    udi4 : inout std_logic;
    udi5 : inout std_logic;
    udi6 : inout std_logic;
    udi7 : inout std_logic;
    udi8 : inout std_logic;
    udi9 : inout std_logic;
    \udo 0\ : out std_logic;
    \udo 1\ : out std_logic;
    \udo 10\ : out std_logic;
    \udo 11\ : out std_logic;
    \udo 12\ : out std_logic;
    \udo 13\ : out std_logic;
    \udo 14\ : out std_logic;
    \udo 15\ : out std_logic;
    \udo 2\ : out std_logic;
    \udo 3\ : out std_logic;
    \udo 4\ : out std_logic;
    \udo 5\ : out std_logic;
    \udo 6\ : out std_logic;
    \udo 7\ : out std_logic;
    \udo 8\ : out std_logic;
    \udo 9\ : out std_logic;
    writeok : inout std_logic
  );
end entity;
