library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn74244_tb is
end sn74244_tb;

architecture testbench of sn74244_tb is

begin

--  uut : sn74244 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
