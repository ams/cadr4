library ieee;
use ieee.std_logic_1164.all;

entity icmem_olord1 is
  port (
    \-boot\         : in     std_logic;
    \-clock reset a\ : in     std_logic;
    \-errhalt\      : in     std_logic;
    \-ldclk\        : in     std_logic;
    \-ldmode\       : in     std_logic;
    \-ldopc\        : in     std_logic;
    \-reset\        : in     std_logic;
    \-stc32\        : in     std_logic;
    \-tpr60\        : in     std_logic;
    \-wait\         : in     std_logic;
    mclk5a          : in     std_logic;
    spy0            : in     std_logic;
    spy1            : in     std_logic;
    spy2            : in     std_logic;
    spy3            : in     std_logic;
    spy4            : in     std_logic;
    spy5            : in     std_logic;
    statstop        : in     std_logic;
    \-idebug\       : out    std_logic;
    \-ldstat\       : out    std_logic;
    \-lpc.hold\     : out    std_logic;
    \-machrun\      : out    std_logic;
    \-machruna\     : out    std_logic;
    \-nop11\        : out    std_logic;
    \-opcclk\       : out    std_logic;
    \-opcinh\       : out    std_logic;
    \-run\          : out    std_logic;
    \-ssdone\       : out    std_logic;
    \-stathalt\     : out    std_logic;
    \-step\         : out    std_logic;
    \lpc.hold\      : out    std_logic;
    \stat.ovf\      : out    std_logic;
    errstop         : out    std_logic;
    idebug          : out    std_logic;
    ldstat          : out    std_logic;
    machrun         : out    std_logic;
    nop11           : out    std_logic;
    opcclk          : out    std_logic;
    opcinh          : out    std_logic;
    promdisable     : out    std_logic;
    promdisabled    : out    std_logic;
    run             : out    std_logic;
    speed0          : out    std_logic;
    speed0a         : out    std_logic;
    speed1          : out    std_logic;
    speed1a         : out    std_logic;
    speedclk        : out    std_logic;
    srun            : out    std_logic;
    ssdone          : out    std_logic;
    sspeed0         : out    std_logic;
    sspeed1         : out    std_logic;
    sstep           : out    std_logic;
    stathenb        : out    std_logic;
    step            : out    std_logic;
    trapenb         : out    std_logic
  );
end entity;
