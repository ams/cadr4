-- CADR1_LMDATA
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_lmdata is
  port (
    \-lmbus enb\ : inout std_logic;
    \bus 0\ : inout std_logic;
    \bus 1\ : inout std_logic;
    \bus 10\ : inout std_logic;
    \bus 11\ : inout std_logic;
    \bus 12\ : inout std_logic;
    \bus 13\ : inout std_logic;
    \bus 14\ : inout std_logic;
    \bus 15\ : inout std_logic;
    \bus 16\ : inout std_logic;
    \bus 17\ : inout std_logic;
    \bus 18\ : inout std_logic;
    \bus 19\ : inout std_logic;
    \bus 2\ : inout std_logic;
    \bus 20\ : inout std_logic;
    \bus 21\ : inout std_logic;
    \bus 22\ : inout std_logic;
    \bus 23\ : inout std_logic;
    \bus 24\ : inout std_logic;
    \bus 25\ : inout std_logic;
    \bus 26\ : inout std_logic;
    \bus 27\ : inout std_logic;
    \bus 28\ : inout std_logic;
    \bus 29\ : inout std_logic;
    \bus 3\ : inout std_logic;
    \bus 30\ : inout std_logic;
    \bus 31\ : inout std_logic;
    \bus 4\ : inout std_logic;
    \bus 5\ : inout std_logic;
    \bus 6\ : inout std_logic;
    \bus 7\ : inout std_logic;
    \bus 8\ : inout std_logic;
    \bus 9\ : inout std_logic;
    \bus _ lm\ : inout std_logic;
    \mem 0\ : inout std_logic;
    \mem 1\ : inout std_logic;
    \mem 10\ : inout std_logic;
    \mem 11\ : inout std_logic;
    \mem 12\ : inout std_logic;
    \mem 13\ : inout std_logic;
    \mem 14\ : inout std_logic;
    \mem 15\ : inout std_logic;
    \mem 16\ : inout std_logic;
    \mem 17\ : inout std_logic;
    \mem 18\ : inout std_logic;
    \mem 19\ : inout std_logic;
    \mem 2\ : inout std_logic;
    \mem 20\ : inout std_logic;
    \mem 21\ : inout std_logic;
    \mem 22\ : inout std_logic;
    \mem 23\ : inout std_logic;
    \mem 24\ : inout std_logic;
    \mem 25\ : inout std_logic;
    \mem 26\ : inout std_logic;
    \mem 27\ : inout std_logic;
    \mem 28\ : inout std_logic;
    \mem 29\ : inout std_logic;
    \mem 3\ : inout std_logic;
    \mem 30\ : inout std_logic;
    \mem 31\ : inout std_logic;
    \mem 4\ : inout std_logic;
    \mem 5\ : inout std_logic;
    \mem 6\ : inout std_logic;
    \mem 7\ : inout std_logic;
    \mem 8\ : inout std_logic;
    \mem 9\ : inout std_logic;
    \mempar from lm\ : inout std_logic
  );
end entity;
