library ieee;
use ieee.std_logic_1164.all;

entity cadr_spcpar is
  port (
    spc0            : in     std_logic;
    spc1            : in     std_logic;
    spc10           : in     std_logic;
    spc11           : in     std_logic;
    spc12           : in     std_logic;
    spc13           : in     std_logic;
    spc14           : in     std_logic;
    spc15           : in     std_logic;
    spc16           : in     std_logic;
    spc17           : in     std_logic;
    spc18           : in     std_logic;
    spc2            : in     std_logic;
    spc3            : in     std_logic;
    spc4            : in     std_logic;
    spc5            : in     std_logic;
    spc6            : in     std_logic;
    spc7            : in     std_logic;
    spc8            : in     std_logic;
    spc9            : in     std_logic;
    spcpar          : in     std_logic;
    spcw0           : in     std_logic;
    spcw1           : in     std_logic;
    spcw10          : in     std_logic;
    spcw11          : in     std_logic;
    spcw12          : in     std_logic;
    spcw13          : in     std_logic;
    spcw14          : in     std_logic;
    spcw15          : in     std_logic;
    spcw16          : in     std_logic;
    spcw17          : in     std_logic;
    spcw18          : in     std_logic;
    spcw2           : in     std_logic;
    spcw3           : in     std_logic;
    spcw4           : in     std_logic;
    spcw5           : in     std_logic;
    spcw6           : in     std_logic;
    spcw7           : in     std_logic;
    spcw8           : in     std_logic;
    spcw9           : in     std_logic;
    \-spcwparl\     : out    std_logic;
    spcparh         : out    std_logic;
    spcparok        : out    std_logic;
    spcwpar         : out    std_logic;
    spcwparh        : out    std_logic
  );
end entity;
