-- Synchronous 4-Bit Up/Down Binary Counter

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Datasheet: Texas Instruments SN74LS169B Synchronous 4-Bit Up/Down Binary Counters, PDIP (N) Package
-- URL: https://www.ti.com/lit/gpn/SN74LS169B

entity sn74169 is
  port (
    co_n : out std_logic;
    i3   : in  std_logic;
    i2   : in  std_logic;
    i1   : in  std_logic;
    i0   : in  std_logic;

    o3      : out std_logic; -- Pin 11 (Output D)
    o2      : out std_logic; -- Pin 12 (Output C)
    o1      : out std_logic; -- Pin 13 (Output B)
    o0      : out std_logic; -- Pin 14 (Output A)

    enb_t_n : in std_logic; -- Pin 10 (Count Enable Trickle Input Active Low)
    enb_p_n : in std_logic; -- Pin 7 (Count Enable Parallel Input Active Low)
    load_n  : in std_logic; -- Pin 9 (Parallel Enable Input Active Low)
    up_dn   : in std_logic; -- Pin 1 (Up/Down Control Input)
    clk     : in std_logic -- Pin 2 (Clock Input)
    );
end;

architecture ttl of sn74169 is
  signal cnt : unsigned(3 downto 0);    -- internal 4-bit register
begin
  ------------------------------------------------------------------
  -- synchronous logic
  ------------------------------------------------------------------
  process(clk)
    variable load_val : unsigned(3 downto 0);
  begin
    if rising_edge(clk) then
      -- synchronous parallel load has top priority
      if load_n = '0' then
        load_val := unsigned'(i3 & i2 & i1 & i0);
        cnt      <= load_val;

      -- otherwise count when both enables are asserted (low)
      elsif (enb_t_n = '0' and enb_p_n = '0') then
        if up_dn = '1' then
          cnt <= cnt + 1;               -- up-count (wraps 15→0)
        else
          cnt <= cnt - 1;               -- down-count (wraps 0→15)
        end if;
      end if;
    -- if enables are not both low, the register simply holds
    end if;
  end process;

  ------------------------------------------------------------------
  -- pin drivers
  ------------------------------------------------------------------
  o3 <= cnt(3);
  o2 <= cnt(2);
  o1 <= cnt(1);
  o0 <= cnt(0);

  -- terminal count / ripple-carry (active-low)
  -- Terminal count occurs when:
  -- 1. Both enables are active (low)
  -- 2. Either:
  --    a. Loading terminal count value (15 for up-count, 0 for down-count)
  --    b. Counter is at terminal count (15 for up-count, 0 for down-count)
  process(all)
    variable at_terminal_count : boolean;
    variable loading_terminal_count : boolean;
  begin
    -- Check if counter is at terminal count
    if up_dn = '1' then
      at_terminal_count := (cnt = to_unsigned(15, 4));  -- up-count terminal
    else
      at_terminal_count := (cnt = to_unsigned(0, 4));   -- down-count terminal
    end if;
    
    -- Check if loading a terminal count value
    if load_n = '0' then
      if up_dn = '1' then
        loading_terminal_count := (unsigned(i3 & i2 & i1 & i0) = to_unsigned(15, 4));
      else
        loading_terminal_count := (unsigned(i3 & i2 & i1 & i0) = to_unsigned(0, 4));
      end if;
    else
      loading_terminal_count := false;
    end if;
    
    -- Generate carry-out (active low)
    if (enb_t_n = '0' and enb_p_n = '0') and (at_terminal_count or loading_terminal_count) then
      co_n <= '0';  -- Active low terminal count
    else
      co_n <= '1';  -- Not at terminal count
    end if;
  end process;
end architecture;
