library ieee;
use ieee.std_logic_1164.all;

entity cadr_vmas is
  port (
    \-md10\         : in     std_logic;
    \-md11\         : in     std_logic;
    \-md12\         : in     std_logic;
    \-md13\         : in     std_logic;
    \-md14\         : in     std_logic;
    \-md15\         : in     std_logic;
    \-md16\         : in     std_logic;
    \-md17\         : in     std_logic;
    \-md18\         : in     std_logic;
    \-md19\         : in     std_logic;
    \-md20\         : in     std_logic;
    \-md21\         : in     std_logic;
    \-md22\         : in     std_logic;
    \-md23\         : in     std_logic;
    \-md8\          : in     std_logic;
    \-md9\          : in     std_logic;
    \-memstart\     : in     std_logic;
    \-vma10\        : in     std_logic;
    \-vma11\        : in     std_logic;
    \-vma12\        : in     std_logic;
    \-vma13\        : in     std_logic;
    \-vma14\        : in     std_logic;
    \-vma15\        : in     std_logic;
    \-vma16\        : in     std_logic;
    \-vma17\        : in     std_logic;
    \-vma18\        : in     std_logic;
    \-vma19\        : in     std_logic;
    \-vma20\        : in     std_logic;
    \-vma21\        : in     std_logic;
    \-vma22\        : in     std_logic;
    \-vma23\        : in     std_logic;
    \-vma8\         : in     std_logic;
    \-vma9\         : in     std_logic;
    lc10            : in     std_logic;
    lc11            : in     std_logic;
    lc12            : in     std_logic;
    lc13            : in     std_logic;
    lc14            : in     std_logic;
    lc15            : in     std_logic;
    lc16            : in     std_logic;
    lc17            : in     std_logic;
    lc18            : in     std_logic;
    lc19            : in     std_logic;
    lc2             : in     std_logic;
    lc20            : in     std_logic;
    lc21            : in     std_logic;
    lc22            : in     std_logic;
    lc23            : in     std_logic;
    lc24            : in     std_logic;
    lc25            : in     std_logic;
    lc3             : in     std_logic;
    lc4             : in     std_logic;
    lc5             : in     std_logic;
    lc6             : in     std_logic;
    lc7             : in     std_logic;
    lc8             : in     std_logic;
    lc9             : in     std_logic;
    ob0             : in     std_logic;
    ob1             : in     std_logic;
    ob10            : in     std_logic;
    ob11            : in     std_logic;
    ob12            : in     std_logic;
    ob13            : in     std_logic;
    ob14            : in     std_logic;
    ob15            : in     std_logic;
    ob16            : in     std_logic;
    ob17            : in     std_logic;
    ob18            : in     std_logic;
    ob19            : in     std_logic;
    ob2             : in     std_logic;
    ob20            : in     std_logic;
    ob21            : in     std_logic;
    ob22            : in     std_logic;
    ob23            : in     std_logic;
    ob24            : in     std_logic;
    ob25            : in     std_logic;
    ob26            : in     std_logic;
    ob27            : in     std_logic;
    ob28            : in     std_logic;
    ob29            : in     std_logic;
    ob3             : in     std_logic;
    ob30            : in     std_logic;
    ob31            : in     std_logic;
    ob4             : in     std_logic;
    ob5             : in     std_logic;
    ob6             : in     std_logic;
    ob7             : in     std_logic;
    ob8             : in     std_logic;
    ob9             : in     std_logic;
    vmasela         : in     std_logic;
    vmaselb         : in     std_logic;
    \-vmas0\        : out    std_logic;
    \-vmas10\       : out    std_logic;
    \-vmas11\       : out    std_logic;
    \-vmas12\       : out    std_logic;
    \-vmas13\       : out    std_logic;
    \-vmas14\       : out    std_logic;
    \-vmas15\       : out    std_logic;
    \-vmas16\       : out    std_logic;
    \-vmas17\       : out    std_logic;
    \-vmas18\       : out    std_logic;
    \-vmas19\       : out    std_logic;
    \-vmas1\        : out    std_logic;
    \-vmas20\       : out    std_logic;
    \-vmas21\       : out    std_logic;
    \-vmas22\       : out    std_logic;
    \-vmas23\       : out    std_logic;
    \-vmas24\       : out    std_logic;
    \-vmas25\       : out    std_logic;
    \-vmas26\       : out    std_logic;
    \-vmas27\       : out    std_logic;
    \-vmas28\       : out    std_logic;
    \-vmas29\       : out    std_logic;
    \-vmas2\        : out    std_logic;
    \-vmas30\       : out    std_logic;
    \-vmas31\       : out    std_logic;
    \-vmas3\        : out    std_logic;
    \-vmas4\        : out    std_logic;
    \-vmas5\        : out    std_logic;
    \-vmas6\        : out    std_logic;
    \-vmas7\        : out    std_logic;
    \-vmas8\        : out    std_logic;
    \-vmas9\        : out    std_logic;
    mapi10          : out    std_logic;
    mapi11          : out    std_logic;
    mapi12          : out    std_logic;
    mapi13          : out    std_logic;
    mapi14          : out    std_logic;
    mapi15          : out    std_logic;
    mapi16          : out    std_logic;
    mapi17          : out    std_logic;
    mapi18          : out    std_logic;
    mapi19          : out    std_logic;
    mapi20          : out    std_logic;
    mapi21          : out    std_logic;
    mapi22          : out    std_logic;
    mapi23          : out    std_logic;
    mapi8           : out    std_logic;
    mapi9           : out    std_logic
  );
end entity;
