library ieee;
use ieee.std_logic_1164.all;

package busint_book is
end package;
