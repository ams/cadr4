library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn7437_tb is
end sn7437_tb;

architecture testbench of sn7437_tb is

begin

--  uut : sn7437 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
