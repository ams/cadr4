library ieee;
use ieee.std_logic_1164.all;

entity cadr_amem1 is
  port (
    \-aadr0a\       : in     std_logic;
    \-aadr1a\       : in     std_logic;
    \-aadr2a\       : in     std_logic;
    \-aadr3a\       : in     std_logic;
    \-aadr4a\       : in     std_logic;
    \-aadr5a\       : in     std_logic;
    \-aadr6a\       : in     std_logic;
    \-aadr7a\       : in     std_logic;
    \-aadr8a\       : in     std_logic;
    \-aadr9a\       : in     std_logic;
    \-awpb\         : in     std_logic;
    \-awpc\         : in     std_logic;
    l0              : in     std_logic;
    l1              : in     std_logic;
    l10             : in     std_logic;
    l11             : in     std_logic;
    l12             : in     std_logic;
    l13             : in     std_logic;
    l14             : in     std_logic;
    l15             : in     std_logic;
    l2              : in     std_logic;
    l3              : in     std_logic;
    l4              : in     std_logic;
    l5              : in     std_logic;
    l6              : in     std_logic;
    l7              : in     std_logic;
    l8              : in     std_logic;
    l9              : in     std_logic;
    amem0           : out    std_logic;
    amem1           : out    std_logic;
    amem10          : out    std_logic;
    amem11          : out    std_logic;
    amem12          : out    std_logic;
    amem13          : out    std_logic;
    amem14          : out    std_logic;
    amem15          : out    std_logic;
    amem2           : out    std_logic;
    amem3           : out    std_logic;
    amem4           : out    std_logic;
    amem5           : out    std_logic;
    amem6           : out    std_logic;
    amem7           : out    std_logic;
    amem8           : out    std_logic;
    amem9           : out    std_logic
  );
end entity cadr_amem1;
