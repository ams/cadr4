library ieee;
use ieee.std_logic_1164.all;

entity busint_rbuf is
  port (
    \-bus>ub\       : in     std_logic;
    \-rbufwe\       : in     std_logic;
    \-ub read buffer\ : in     std_logic;
    \-ubpn0b\       : in     std_logic;
    \-ubpn1b\       : in     std_logic;
    \-ubpn2b\       : in     std_logic;
    \-ubpn3b\       : in     std_logic;
    bus0            : in     std_logic;
    bus1            : in     std_logic;
    bus10           : in     std_logic;
    bus11           : in     std_logic;
    bus12           : in     std_logic;
    bus13           : in     std_logic;
    bus14           : in     std_logic;
    bus15           : in     std_logic;
    bus16           : in     std_logic;
    bus17           : in     std_logic;
    bus18           : in     std_logic;
    bus19           : in     std_logic;
    bus2            : in     std_logic;
    bus20           : in     std_logic;
    bus21           : in     std_logic;
    bus22           : in     std_logic;
    bus23           : in     std_logic;
    bus24           : in     std_logic;
    bus25           : in     std_logic;
    bus26           : in     std_logic;
    bus27           : in     std_logic;
    bus28           : in     std_logic;
    bus29           : in     std_logic;
    bus3            : in     std_logic;
    bus30           : in     std_logic;
    bus31           : in     std_logic;
    bus4            : in     std_logic;
    bus5            : in     std_logic;
    bus6            : in     std_logic;
    bus7            : in     std_logic;
    bus8            : in     std_logic;
    bus9            : in     std_logic;
    rbuf16          : out    std_logic;
    rbuf17          : out    std_logic;
    rbuf18          : out    std_logic;
    rbuf19          : out    std_logic;
    rbuf20          : out    std_logic;
    rbuf21          : out    std_logic;
    rbuf22          : out    std_logic;
    rbuf23          : out    std_logic;
    rbuf24          : out    std_logic;
    rbuf25          : out    std_logic;
    rbuf26          : out    std_logic;
    rbuf27          : out    std_logic;
    rbuf28          : out    std_logic;
    rbuf29          : out    std_logic;
    rbuf30          : out    std_logic;
    rbuf31          : out    std_logic;
    udo0            : out    std_logic;
    udo1            : out    std_logic;
    udo10           : out    std_logic;
    udo11           : out    std_logic;
    udo12           : out    std_logic;
    udo13           : out    std_logic;
    udo14           : out    std_logic;
    udo15           : out    std_logic;
    udo2            : out    std_logic;
    udo3            : out    std_logic;
    udo4            : out    std_logic;
    udo5            : out    std_logic;
    udo6            : out    std_logic;
    udo7            : out    std_logic;
    udo8            : out    std_logic;
    udo9            : out    std_logic
  );
end entity busint_rbuf;
