library ieee;
use ieee.std_logic_1164.all;

entity md is
  port (
    \-mddrive\  : out std_logic;
    \-md31\     : out std_logic;
    mf24        : out std_logic;
    \-md30\     : out std_logic;
    mf25        : out std_logic;
    \-md29\     : out std_logic;
    mf26        : out std_logic;
    \-md28\     : out std_logic;
    mf27        : out std_logic;
    \-md27\     : out std_logic;
    mf28        : out std_logic;
    \-md26\     : out std_logic;
    mf29        : out std_logic;
    \-md25\     : out std_logic;
    mf30        : out std_logic;
    \-md24\     : out std_logic;
    mf31        : out std_logic;
    \-md23\     : out std_logic;
    mf16        : out std_logic;
    \-md22\     : out std_logic;
    mf17        : out std_logic;
    \-md21\     : out std_logic;
    mf18        : out std_logic;
    \-md20\     : out std_logic;
    mf19        : out std_logic;
    \-md19\     : out std_logic;
    mf20        : out std_logic;
    \-md18\     : out std_logic;
    mf21        : out std_logic;
    \-md17\     : out std_logic;
    mf22        : out std_logic;
    \-md16\     : out std_logic;
    mf23        : out std_logic;
    \-md7\      : out std_logic;
    mf0         : out std_logic;
    \-md6\      : out std_logic;
    mf1         : out std_logic;
    \-md5\      : out std_logic;
    mf2         : out std_logic;
    \-md4\      : out std_logic;
    mf3         : out std_logic;
    \-md3\      : out std_logic;
    mf4         : out std_logic;
    \-md2\      : out std_logic;
    mf5         : out std_logic;
    \-md1\      : out std_logic;
    mf6         : out std_logic;
    \-md0\      : out std_logic;
    mf7         : out std_logic;
    srcmd       : out std_logic;
    tse2        : in  std_logic;
    \-md15\     : out std_logic;
    mf8         : out std_logic;
    \-md14\     : out std_logic;
    mf9         : out std_logic;
    \-md13\     : out std_logic;
    mf10        : out std_logic;
    \-md12\     : out std_logic;
    mf11        : out std_logic;
    \-md11\     : out std_logic;
    mf12        : out std_logic;
    \-md10\     : out std_logic;
    mf13        : out std_logic;
    \-md9\      : out std_logic;
    mf14        : out std_logic;
    \-md8\      : out std_logic;
    mf15        : out std_logic;
    gnd         : in  std_logic;
    \-mds31\    : in  std_logic;
    \-mds30\    : in  std_logic;
    \-mds29\    : in  std_logic;
    \-mds28\    : in  std_logic;
    mdclk       : out std_logic;
    \-mds27\    : in  std_logic;
    \-mds26\    : in  std_logic;
    \-mds25\    : in  std_logic;
    \-mds24\    : in  std_logic;
    \-mds7\     : in  std_logic;
    \-mds6\     : in  std_logic;
    \-mds5\     : in  std_logic;
    \-mds4\     : in  std_logic;
    \-mds3\     : in  std_logic;
    \-mds2\     : in  std_logic;
    \-mds1\     : in  std_logic;
    \-mds0\     : in  std_logic;
    \-mds23\    : in  std_logic;
    \-mds22\    : in  std_logic;
    \-mds21\    : in  std_logic;
    \-mds20\    : in  std_logic;
    \-mds19\    : in  std_logic;
    \-mds18\    : in  std_logic;
    \-mds17\    : in  std_logic;
    \-mds16\    : in  std_logic;
    destmdr     : out std_logic;
    \-clk2c\    : in  std_logic;
    loadmd      : out std_logic;
    \-loadmd\   : in  std_logic;
    \-destmdr\  : in  std_logic;
    \-mds15\    : in  std_logic;
    \-mds14\    : in  std_logic;
    \-mds13\    : in  std_logic;
    \-mds12\    : in  std_logic;
    \-mds11\    : in  std_logic;
    \-mds10\    : in  std_logic;
    \-mds9\     : in  std_logic;
    \-mds8\     : in  std_logic;
    mdgetspar   : out std_logic;
    \-ignpar\   : in  std_logic;
    mdhaspar    : out std_logic;
    \mempar_in\ : in  std_logic;
    mdpar       : out std_logic;
    \-srcmd\    : in  std_logic);
end;
