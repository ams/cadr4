library ieee;
use ieee.std_logic_1164.all;

entity cadr_pdlctl is
  port (
    \-reset\      : in  std_logic;
    pdlwrited     : out std_logic;
    \-pdlwrited\  : out std_logic;
    pdlwrite      : out std_logic;
    \-destpdl(x)\ : in  std_logic;
    pwidx         : out std_logic;
    \-pwidx\      : out std_logic;
    clk4f         : in  std_logic;
    imodd         : out std_logic;
    \-imodd\      : out std_logic;
    imod          : in  std_logic;
    \-destspc\    : in  std_logic;
    \-destspcd\   : out std_logic;
    \-pdlpb\      : out std_logic;
    pdlptr0       : in  std_logic;
    pdlidx0       : in  std_logic;
    \-pdla0b\     : out std_logic;
    pdlptr1       : in  std_logic;
    pdlidx1       : in  std_logic;
    \-pdla1b\     : out std_logic;
    \-pdla2b\     : out std_logic;
    pdlidx2       : in  std_logic;
    pdlptr2       : in  std_logic;
    \-pdla3b\     : out std_logic;
    pdlidx3       : in  std_logic;
    pdlptr3       : in  std_logic;
    gnd           : in  std_logic;
    \-pdlpa\      : out std_logic;
    pdlptr8       : in  std_logic;
    pdlidx8       : in  std_logic;
    \-pdla8b\     : out std_logic;
    pdlptr9       : in  std_logic;
    pdlidx9       : in  std_logic;
    \-pdla9b\     : out std_logic;
    \-pdla0a\     : out std_logic;
    \-pdla1a\     : out std_logic;
    \-pdla2a\     : out std_logic;
    \-pdla3a\     : out std_logic;
    \-pdla4a\     : out std_logic;
    pdlidx4       : in  std_logic;
    pdlptr4       : in  std_logic;
    \-pdla5a\     : out std_logic;
    pdlidx5       : in  std_logic;
    pdlptr5       : in  std_logic;
    \-destpdl(p)\ : in  std_logic;
    \-pdlcnt\     : out std_logic;
    clk4b         : in  std_logic;
    ir30          : in  std_logic;
    \-clk4e\      : in  std_logic;
    \-srcpdlpop\  : in  std_logic;
    \-srcpdltop\  : in  std_logic;
    pdlenb        : out std_logic;
    tse4b         : in  std_logic;
    \-pdldrive\   : out std_logic;
    \-destpdltop\ : in  std_logic;
    \-pdla4b\     : out std_logic;
    \-pdla5b\     : out std_logic;
    \-pdla6b\     : out std_logic;
    pdlidx6       : in  std_logic;
    pdlptr6       : in  std_logic;
    \-pdla7b\     : out std_logic;
    pdlidx7       : in  std_logic;
    pdlptr7       : in  std_logic;
    wp4a          : in  std_logic;
    \-pwpa\       : out std_logic;
    \-pwpb\       : out std_logic;
    \-pwpc\       : out std_logic;
    \-pdla6a\     : out std_logic;
    \-pdla7a\     : out std_logic;
    \-pdla8a\     : out std_logic;
    \-pdla9a\     : out std_logic;
    nop           : in  std_logic);
end;
