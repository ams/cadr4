library ieee;
use ieee.std_logic_1164.all;

entity cadr_mds is
  port (
    \-memdrive.a\ : in  std_logic;
    \-md31\       : in  std_logic;
    mem24         : out std_logic;
    \-md30\       : in  std_logic;
    mem25         : out std_logic;
    \-md29\       : in  std_logic;
    mem26         : out std_logic;
    \-md28\       : in  std_logic;
    \-md27\       : in  std_logic;
    mem28         : out std_logic;
    \-md26\       : in  std_logic;
    mem29         : out std_logic;
    \-md25\       : in  std_logic;
    mem30         : out std_logic;
    \-md24\       : in  std_logic;
    mem31         : out std_logic;
    \-memdrive.b\ : in  std_logic;
    \-md7\        : in  std_logic;
    mem0          : out std_logic;
    \-md6\        : in  std_logic;
    mem1          : out std_logic;
    \-md5\        : in  std_logic;
    mem2          : out std_logic;
    \-md4\        : in  std_logic;
    mem3          : out std_logic;
    \-md3\        : in  std_logic;
    mem4          : out std_logic;
    \-md2\        : in  std_logic;
    mem5          : out std_logic;
    \-md1\        : in  std_logic;
    mem6          : out std_logic;
    \-md0\        : in  std_logic;
    mem7          : out std_logic;
    \-md23\       : in  std_logic;
    mem16         : out std_logic;
    \-md22\       : in  std_logic;
    mem17         : out std_logic;
    \-md21\       : in  std_logic;
    mem18         : out std_logic;
    \-md20\       : in  std_logic;
    mem19         : out std_logic;
    \-md19\       : in  std_logic;
    mem20         : out std_logic;
    \-md18\       : in  std_logic;
    mem21         : out std_logic;
    \-md17\       : in  std_logic;
    mem22         : out std_logic;
    \-md16\       : in  std_logic;
    mem23         : out std_logic;
    \-md15\       : in  std_logic;
    mem8          : out std_logic;
    \-md14\       : in  std_logic;
    mem9          : out std_logic;
    \-md13\       : in  std_logic;
    mem10         : out std_logic;
    \-md12\       : in  std_logic;
    mem11         : out std_logic;
    \-md11\       : in  std_logic;
    mem12         : out std_logic;
    \-md10\       : in  std_logic;
    mem13         : out std_logic;
    \-md9\        : in  std_logic;
    mem14         : out std_logic;
    \-md8\        : in  std_logic;
    mem15         : out std_logic;
    mdsela        : in  std_logic;
    ob20          : in  std_logic;
    \-mds20\      : out std_logic;
    ob21          : in  std_logic;
    \-mds21\      : out std_logic;
    \-mds22\      : out std_logic;
    ob22          : in  std_logic;
    \-mds23\      : out std_logic;
    ob23          : in  std_logic;
    gnd           : in  std_logic;
    ob28          : in  std_logic;
    \-mds28\      : out std_logic;
    ob29          : in  std_logic;
    \-mds29\      : out std_logic;
    \-mds30\      : out std_logic;
    ob30          : in  std_logic;
    \-mds31\      : out std_logic;
    ob31          : in  std_logic;
    mdparodd      : in  std_logic;
    \mempar out\  : out std_logic;
    hi11          : in  std_logic;
    mdselb        : in  std_logic;
    ob12          : in  std_logic;
    \-mds12\      : out std_logic;
    ob13          : in  std_logic;
    \-mds13\      : out std_logic;
    \-mds14\      : out std_logic;
    ob14          : in  std_logic;
    \-mds15\      : out std_logic;
    ob15          : in  std_logic;
    ob16          : in  std_logic;
    \-mds16\      : out std_logic;
    ob17          : in  std_logic;
    \-mds17\      : out std_logic;
    \-mds18\      : out std_logic;
    ob18          : in  std_logic;
    \-mds19\      : out std_logic;
    ob19          : in  std_logic;
    ob8           : in  std_logic;
    \-mds8\       : out std_logic;
    ob9           : in  std_logic;
    \-mds9\       : out std_logic;
    \-mds10\      : out std_logic;
    ob10          : in  std_logic;
    \-mds11\      : out std_logic;
    ob11          : in  std_logic;
    ob0           : in  std_logic;
    \-mds0\       : out std_logic;
    ob1           : in  std_logic;
    \-mds1\       : out std_logic;
    \-mds2\       : out std_logic;
    ob2           : in  std_logic;
    \-mds3\       : out std_logic;
    ob3           : in  std_logic;
    ob4           : in  std_logic;
    \-mds4\       : out std_logic;
    ob5           : in  std_logic;
    \-mds5\       : out std_logic;
    \-mds6\       : out std_logic;
    ob6           : in  std_logic;
    \-mds7\       : out std_logic;
    ob7           : in  std_logic;
    ob24          : in  std_logic;
    \-mds24\      : out std_logic;
    ob25          : in  std_logic;
    \-mds25\      : out std_logic;
    \-mds26\      : out std_logic;
    ob26          : in  std_logic;
    \-mds27\      : out std_logic;
    ob27          : in  std_logic;
    mem27         : out std_logic
    );
end;
