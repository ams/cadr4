library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_mlatch is
  port (
    \-mpassm\  : in  std_logic;
    m23        : out std_logic;
    mmem23     : in  std_logic;
    mmem22     : out std_logic;
    m22        : out std_logic;
    m21        : out std_logic;
    mmem21     : in  std_logic;
    mmem20     : out std_logic;
    m20        : out std_logic;
    clk4a      : in  std_logic;
    m19        : out std_logic;
    mmem19     : in  std_logic;
    mmem18     : out std_logic;
    m18        : out std_logic;
    m17        : out std_logic;
    mmem17     : in  std_logic;
    mmem16     : out std_logic;
    m16        : out std_logic;
    m15        : out std_logic;
    mmem15     : in  std_logic;
    mmem14     : out std_logic;
    m14        : out std_logic;
    m13        : out std_logic;
    mmem13     : in  std_logic;
    mmem12     : out std_logic;
    m12        : out std_logic;
    m11        : out std_logic;
    mmem11     : in  std_logic;
    mmem10     : out std_logic;
    m10        : out std_logic;
    m9         : out std_logic;
    mmem9      : in  std_logic;
    mmem8      : out std_logic;
    m8         : out std_logic;
    m7         : out std_logic;
    mmem7      : in  std_logic;
    mmem6      : out std_logic;
    m6         : out std_logic;
    m5         : out std_logic;
    mmem5      : in  std_logic;
    mmem4      : out std_logic;
    m4         : out std_logic;
    m3         : out std_logic;
    mmem3      : in  std_logic;
    mmem2      : in  std_logic;
    m2         : out std_logic;
    m1         : out std_logic;
    mmem1      : out std_logic;
    mmem0      : out std_logic;
    m0         : out std_logic;
    \-mpassl\  : in  std_logic;
    l15        : in  std_logic;
    mf8        : out std_logic;
    l14        : in  std_logic;
    mf9        : out std_logic;
    l13        : in  std_logic;
    mf10       : out std_logic;
    l12        : in  std_logic;
    mf11       : out std_logic;
    l11        : in  std_logic;
    mf12       : out std_logic;
    l10        : in  std_logic;
    mf13       : out std_logic;
    l9         : in  std_logic;
    mf14       : out std_logic;
    l8         : in  std_logic;
    mf15       : out std_logic;
    mpassl     : in  std_logic;
    l7         : in  std_logic;
    mf0        : out std_logic;
    l6         : in  std_logic;
    mf1        : out std_logic;
    l5         : in  std_logic;
    mf2        : out std_logic;
    l4         : in  std_logic;
    mf3        : out std_logic;
    l3         : in  std_logic;
    mf4        : out std_logic;
    l2         : in  std_logic;
    mf5        : out std_logic;
    l1         : in  std_logic;
    mf6        : out std_logic;
    l0         : in  std_logic;
    mf7        : out std_logic;
    mmemparity : out std_logic;
    mparity    : out std_logic;
    m31        : out std_logic;
    mmem31     : in  std_logic;
    mmem30     : out std_logic;
    m30        : out std_logic;
    m29        : out std_logic;
    mmem29     : in  std_logic;
    mmem28     : out std_logic;
    m28        : out std_logic;
    m27        : out std_logic;
    mmem27     : in  std_logic;
    mmem26     : out std_logic;
    m26        : out std_logic;
    m25        : out std_logic;
    mmem25     : in  std_logic;
    mmem24     : out std_logic;
    m24        : out std_logic;
    l31        : in  std_logic;
    mf24       : out std_logic;
    l30        : in  std_logic;
    mf25       : out std_logic;
    l29        : in  std_logic;
    mf26       : out std_logic;
    l28        : in  std_logic;
    mf27       : out std_logic;
    l27        : in  std_logic;
    mf28       : out std_logic;
    l26        : in  std_logic;
    mf29       : out std_logic;
    l25        : in  std_logic;
    mf30       : out std_logic;
    l24        : in  std_logic;
    mf31       : out std_logic;
    l23        : in  std_logic;
    mf16       : out std_logic;
    l22        : in  std_logic;
    mf17       : out std_logic;
    l21        : in  std_logic;
    mf18       : out std_logic;
    l20        : in  std_logic;
    mf19       : out std_logic;
    l19        : in  std_logic;
    mf20       : out std_logic;
    l18        : in  std_logic;
    mf21       : out std_logic;
    l17        : in  std_logic;
    mf22       : out std_logic;
    l16        : in  std_logic;
    mf23       : out std_logic);
end;

architecture ttl of cadr4_mlatch is
  signal nc294 : std_logic;
  signal nc295 : std_logic;
  signal nc296 : std_logic;
  signal nc297 : std_logic;
  signal nc298 : std_logic;
  signal nc299 : std_logic;
  signal nc300 : std_logic;
  signal nc301 : std_logic;
  signal nc302 : std_logic;
  signal nc303 : std_logic;
  signal nc304 : std_logic;
  signal nc305 : std_logic;
  signal nc306 : std_logic;
  signal nc307 : std_logic;
begin
  mlatch_4a01 : sn74s373 port map(oenb_n => \-mpassm\, o0 => m23, i0 => mmem23, i1 => mmem22, o1 => m22, o2 => m21, i2 => mmem21, i3 => mmem20, o3 => m20, hold_n => clk4a, o4 => m19, i4 => mmem19, i5 => mmem18, o5 => m18, o6 => m17, i6 => mmem17, i7 => mmem16, o7 => m16);
  mlatch_4a03 : sn74s373 port map(oenb_n => \-mpassm\, o0 => m15, i0 => mmem15, i1 => mmem14, o1 => m14, o2 => m13, i2 => mmem13, i3 => mmem12, o3 => m12, hold_n => clk4a, o4 => m11, i4 => mmem11, i5 => mmem10, o5 => m10, o6 => m9, i6 => mmem9, i7 => mmem8, o7 => m8);
  mlatch_4a05 : sn74s373 port map(oenb_n => \-mpassm\, o0 => m7, i0 => mmem7, i1 => mmem6, o1 => m6, o2 => m5, i2 => mmem5, i3 => mmem4, o3 => m4, hold_n => clk4a, o4 => m3, i4 => mmem3, i5 => mmem2, o5 => m2, o6 => m1, i6 => mmem1, i7 => mmem0, o7 => m0);
  mlatch_4a06 : sn74s241 port map(aenb_n => \-mpassl\, ain0 => l15, bout3 => mf8, ain1 => l14, bout2 => mf9, ain2 => l13, bout1 => mf10, ain3 => l12, bout0 => mf11, bin0 => l11, aout3 => mf12, bin1 => l10, aout2 => mf13, bin2 => l9, aout1 => mf14, bin3 => l8, aout0 => mf15, benb => mpassl);
  mlatch_4a08 : sn74s241 port map(aenb_n => \-mpassl\, ain0 => l7, bout3 => mf0, ain1 => l6, bout2 => mf1, ain2 => l5, bout1 => mf2, ain3 => l4, bout0 => mf3, bin0 => l3, aout3 => mf4, bin1 => l2, aout2 => mf5, bin2 => l1, aout1 => mf6, bin3 => l0, aout0 => mf7, benb => mpassl);
  mlatch_4b02 : sn74s373 port map(oenb_n => \-mpassm\, o0 => nc294, i0 => nc295, i1 => nc296, o1 => nc297, o2 => nc298, i2 => nc299, i3 => nc300, o3 => nc301, hold_n => clk4a, o4 => nc302, i4 => nc303, i5 => nc304, o5 => nc305, o6 => nc306, i6 => nc307, i7 => mmemparity, o7 => mparity);
  mlatch_4b04 : sn74s373 port map(oenb_n => \-mpassm\, o0 => m31, i0 => mmem31, i1 => mmem30, o1 => m30, o2 => m29, i2 => mmem29, i3 => mmem28, o3 => m28, hold_n => clk4a, o4 => m27, i4 => mmem27, i5 => mmem26, o5 => m26, o6 => m25, i6 => mmem25, i7 => mmem24, o7 => m24);
  mlatch_4b07 : sn74s241 port map(aenb_n => \-mpassl\, ain0 => l31, bout3 => mf24, ain1 => l30, bout2 => mf25, ain2 => l29, bout1 => mf26, ain3 => l28, bout0 => mf27, bin0 => l27, aout3 => mf28, bin1 => l26, aout2 => mf29, bin2 => l25, aout1 => mf30, bin3 => l24, aout0 => mf31, benb => mpassl);
  mlatch_4b09 : sn74s241 port map(aenb_n => \-mpassl\, ain0 => l23, bout3 => mf16, ain1 => l22, bout2 => mf17, ain2 => l21, bout1 => mf18, ain3 => l20, bout0 => mf19, bin0 => l19, aout3 => mf20, bin1 => l18, aout2 => mf21, bin2 => l17, aout1 => mf22, bin3 => l16, aout0 => mf23, benb => mpassl);
end architecture;
