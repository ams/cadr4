library ieee;
use ieee.std_logic_1164.all;

package busint_book is

  component cadr1_buspar is
  port (
      bus0            : in     std_logic;
      bus1            : in     std_logic;
      bus10           : in     std_logic;
      bus11           : in     std_logic;
      bus12           : in     std_logic;
      bus13           : in     std_logic;
      bus14           : in     std_logic;
      bus15           : in     std_logic;
      bus16           : in     std_logic;
      bus17           : in     std_logic;
      bus18           : in     std_logic;
      bus19           : in     std_logic;
      bus2            : in     std_logic;
      bus20           : in     std_logic;
      bus21           : in     std_logic;
      bus22           : in     std_logic;
      bus23           : in     std_logic;
      bus24           : in     std_logic;
      bus25           : in     std_logic;
      bus26           : in     std_logic;
      bus27           : in     std_logic;
      bus28           : in     std_logic;
      bus29           : in     std_logic;
      bus3            : in     std_logic;
      bus30           : in     std_logic;
      bus31           : in     std_logic;
      bus4            : in     std_logic;
      bus5            : in     std_logic;
      bus6            : in     std_logic;
      bus7            : in     std_logic;
      bus8            : in     std_logic;
      bus9            : in     std_logic;
      \bus 0-11 par odd\ : inout  std_logic;
      \bus 12-23 par odd\ : inout  std_logic;
      \bus par even\  : out    std_logic;
      \bus par odd\   : out    std_logic
    );
  end component;

  component cadr1_bussel is
  port (
      \-ub16>bus\     : in     std_logic;
      \-ub32>bus\     : in     std_logic;
      udi0            : in     std_logic;
      udi1            : in     std_logic;
      udi10           : in     std_logic;
      udi11           : in     std_logic;
      udi12           : in     std_logic;
      udi13           : in     std_logic;
      udi14           : in     std_logic;
      udi15           : in     std_logic;
      udi2            : in     std_logic;
      udi3            : in     std_logic;
      udi4            : in     std_logic;
      udi5            : in     std_logic;
      udi6            : in     std_logic;
      udi7            : in     std_logic;
      udi8            : in     std_logic;
      udi9            : in     std_logic;
      wbuf0           : in     std_logic;
      wbuf1           : in     std_logic;
      wbuf10          : in     std_logic;
      wbuf11          : in     std_logic;
      wbuf12          : in     std_logic;
      wbuf13          : in     std_logic;
      wbuf14          : in     std_logic;
      wbuf15          : in     std_logic;
      wbuf2           : in     std_logic;
      wbuf3           : in     std_logic;
      wbuf4           : in     std_logic;
      wbuf5           : in     std_logic;
      wbuf6           : in     std_logic;
      wbuf7           : in     std_logic;
      wbuf8           : in     std_logic;
      wbuf9           : in     std_logic;
      bus0            : out    std_logic;
      bus1            : out    std_logic;
      bus10           : out    std_logic;
      bus11           : out    std_logic;
      bus12           : out    std_logic;
      bus13           : out    std_logic;
      bus14           : out    std_logic;
      bus15           : out    std_logic;
      bus16           : out    std_logic;
      bus17           : out    std_logic;
      bus18           : out    std_logic;
      bus19           : out    std_logic;
      bus2            : out    std_logic;
      bus20           : out    std_logic;
      bus21           : out    std_logic;
      bus22           : out    std_logic;
      bus23           : out    std_logic;
      bus24           : out    std_logic;
      bus25           : out    std_logic;
      bus26           : out    std_logic;
      bus27           : out    std_logic;
      bus28           : out    std_logic;
      bus29           : out    std_logic;
      bus3            : out    std_logic;
      bus30           : out    std_logic;
      bus31           : out    std_logic;
      bus4            : out    std_logic;
      bus5            : out    std_logic;
      bus6            : out    std_logic;
      bus7            : out    std_logic;
      bus8            : out    std_logic;
      bus9            : out    std_logic
    );
  end component;

  component cadr1_clm is
  port (
      \-mclk7\        : inout  std_logic;
      \-memrq\        : inout  std_logic;
      \-xbus power reset\ : inout  std_logic;
      \hi 15-30\      : inout  std_logic;
      clk0            : inout  std_logic;
      wrcyc           : inout  std_logic;
      \-clk\          : out    std_logic
    );
  end component;

  component cadr1_datctl is
  port (
      \-dbub master\  : in     std_logic;
      \-select debug\ : in     std_logic;
      \-select spy\   : in     std_logic;
      \-ub write buffer\ : in     std_logic;
      \-write through\ : in     std_logic;
      \c1 in\         : in     std_logic;
      \dbub master\   : in     std_logic;
      \debug in wr\   : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \int busy\      : in     std_logic;
      \lmub grant\    : in     std_logic;
      \lmub master\   : in     std_logic;
      \lmx grant a\   : in     std_logic;
      \lmx grant\     : in     std_logic;
      \msyn in\       : in     std_logic;
      \select debug\  : in     std_logic;
      \select page\   : in     std_logic;
      \ub reg cyc t0\ : in     std_logic;
      \ub reg cyc t150\ : in     std_logic;
      \ub reg write pulse\ : in     std_logic;
      \ub17-14=map\   : in     std_logic;
      \ubrd a\        : in     std_logic;
      \ubx grant a\   : in     std_logic;
      \ubx grant\     : in     std_logic;
      lmrd            : in     std_logic;
      lmwr            : in     std_logic;
      ubrd            : in     std_logic;
      ubwr            : in     std_logic;
      wrcyc           : in     std_logic;
      \-ubdrive\      : inout  std_logic;
      \-ubwr\         : inout  std_logic;
      \-xdrive\       : inout  std_logic;
      \write data > ub\ : inout  std_logic;
      \write through\ : inout  std_logic;
      \-bus>ub\       : out    std_logic;
      \-lmadr>ub\     : out    std_logic;
      \-lmadr>xbus\   : out    std_logic;
      \-lmbus enb\    : out    std_logic;
      \-lmrd\         : out    std_logic;
      \-lmwr\         : out    std_logic;
      \-ub16>bus\     : out    std_logic;
      \-ub32>bus\     : out    std_logic;
      \-ubaddr>xbus\  : out    std_logic;
      \-ubadrive\     : out    std_logic;
      \-ubmap > udo\  : out    std_logic;
      \-ubmapwe\      : out    std_logic;
      \-ubrd\         : out    std_logic;
      \-ubwr a\       : out    std_logic;
      \-udi > udo\    : out    std_logic;
      \-wbufwe\       : out    std_logic;
      \-xaddrdrive\   : out    std_logic;
      \-xb>bus\       : out    std_logic;
      \bus > lm\      : out    std_logic;
      xwr             : out    std_logic
    );
  end component;

  component cadr1_dbgin is
  port (
      \-dbub master\  : in     std_logic;
      \-debug reset\  : in     std_logic;
      \-lm power reset\ : in     std_logic;
      \-lm unibus reset\ : in     std_logic;
      \dbub master\   : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \hi 15-30\      : in     std_logic;
      \ssyn t0\       : in     std_logic;
      \unibus init in\ : in     std_logic;
      dbd0            : in     std_logic;
      dbd1            : in     std_logic;
      dbd10           : in     std_logic;
      dbd11           : in     std_logic;
      dbd12           : in     std_logic;
      dbd13           : in     std_logic;
      dbd14           : in     std_logic;
      dbd15           : in     std_logic;
      dbd2            : in     std_logic;
      dbd3            : in     std_logic;
      dbd4            : in     std_logic;
      dbd5            : in     std_logic;
      dbd6            : in     std_logic;
      dbd7            : in     std_logic;
      dbd8            : in     std_logic;
      dbd9            : in     std_logic;
      \-db adr0 clk\  : inout  std_logic;
      \-db adr1 clk\  : inout  std_logic;
      \-db need ub\   : inout  std_logic;
      \-db read status\ : inout  std_logic;
      \-debug in req\ : inout  std_logic;
      \-debugee reset\ : inout  std_logic;
      \-local enable\ : inout  std_logic;
      \debug in a0\   : inout  std_logic;
      \debug in a1\   : inout  std_logic;
      \debug in wr\   : inout  std_logic;
      \debug out ack\ : inout  std_logic;
      \local enable\  : inout  std_logic;
      reset           : inout  std_logic;
      \-busint lm reset\ : out    std_logic;
      \-debug timeout inh\ : out    std_logic;
      \-reset\        : out    std_logic;
      \db need ub\    : out    std_logic;
      \debug ack\     : out    std_logic;
      uao1            : out    std_logic;
      uao10           : out    std_logic;
      uao11           : out    std_logic;
      uao12           : out    std_logic;
      uao13           : out    std_logic;
      uao14           : out    std_logic;
      uao15           : out    std_logic;
      uao16           : out    std_logic;
      uao17           : out    std_logic;
      uao2            : out    std_logic;
      uao3            : out    std_logic;
      uao4            : out    std_logic;
      uao5            : out    std_logic;
      uao6            : out    std_logic;
      uao7            : out    std_logic;
      uao8            : out    std_logic;
      uao9            : out    std_logic
    );
  end component;

  component cadr1_dbgout is
  port (
      \-select debug\ : in     std_logic;
      \dbub master\   : in     std_logic;
      \debug ack\     : in     std_logic;
      \debug in wr\   : in     std_logic;
      \debug out ack\ : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \hi 15-30\      : in     std_logic;
      \select debug dlyd\ : in     std_logic;
      \ud > debug\    : in     std_logic;
      \xbus par in\   : in     std_logic;
      dbd0            : in     std_logic;
      dbd1            : in     std_logic;
      dbd10           : in     std_logic;
      dbd11           : in     std_logic;
      dbd12           : in     std_logic;
      dbd13           : in     std_logic;
      dbd14           : in     std_logic;
      dbd15           : in     std_logic;
      dbd2            : in     std_logic;
      dbd3            : in     std_logic;
      dbd4            : in     std_logic;
      dbd5            : in     std_logic;
      dbd6            : in     std_logic;
      dbd7            : in     std_logic;
      dbd8            : in     std_logic;
      dbd9            : in     std_logic;
      uba1            : in     std_logic;
      uba2            : in     std_logic;
      uba3            : in     std_logic;
      uba4            : in     std_logic;
      ubrd            : in     std_logic;
      ubwr            : in     std_logic;
      udo0            : in     std_logic;
      udo1            : in     std_logic;
      udo10           : in     std_logic;
      udo11           : in     std_logic;
      udo12           : in     std_logic;
      udo13           : in     std_logic;
      udo14           : in     std_logic;
      udo15           : in     std_logic;
      udo2            : in     std_logic;
      udo3            : in     std_logic;
      udo4            : in     std_logic;
      udo5            : in     std_logic;
      udo6            : in     std_logic;
      udo7            : in     std_logic;
      udo8            : in     std_logic;
      udo9            : in     std_logic;
      \-dbd enb\      : inout  std_logic;
      \debug active\  : inout  std_logic;
      \select debug\  : inout  std_logic;
      \-debug > ud\   : out    std_logic;
      \-debug out req\ : out    std_logic;
      \debug in ack\  : out    std_logic;
      \debug out a0\  : out    std_logic;
      \debug out a1\  : out    std_logic;
      \debug out wr\  : out    std_logic;
      \debug ssyn\    : out    std_logic;
      \mempar to lm\  : out    std_logic;
      \spy adr1\      : out    std_logic;
      \spy adr2\      : out    std_logic;
      \spy adr3\      : out    std_logic;
      \spy adr4\      : out    std_logic
    );
  end component;

  component cadr1_diag is
  port (
      \-select spy\   : in     std_logic;
      \ub reg write pulse\ : in     std_logic;
      spy0            : in     std_logic;
      spy1            : in     std_logic;
      spy10           : in     std_logic;
      spy11           : in     std_logic;
      spy12           : in     std_logic;
      spy13           : in     std_logic;
      spy14           : in     std_logic;
      spy15           : in     std_logic;
      spy2            : in     std_logic;
      spy3            : in     std_logic;
      spy4            : in     std_logic;
      spy5            : in     std_logic;
      spy6            : in     std_logic;
      spy7            : in     std_logic;
      spy8            : in     std_logic;
      spy9            : in     std_logic;
      ubrd            : in     std_logic;
      ubwr            : in     std_logic;
      udo0            : in     std_logic;
      udo1            : in     std_logic;
      udo10           : in     std_logic;
      udo11           : in     std_logic;
      udo12           : in     std_logic;
      udo13           : in     std_logic;
      udo14           : in     std_logic;
      udo15           : in     std_logic;
      udo2            : in     std_logic;
      udo3            : in     std_logic;
      udo4            : in     std_logic;
      udo5            : in     std_logic;
      udo6            : in     std_logic;
      udo7            : in     std_logic;
      udo8            : in     std_logic;
      udo9            : in     std_logic;
      \select spy\    : inout  std_logic;
      \-spy read\     : out    std_logic;
      \-spy write\    : out    std_logic
    );
  end component;

  component cadr1_lmadr is
  port (
      \-adr0\         : in     std_logic;
      \-adr10\        : in     std_logic;
      \-adr11\        : in     std_logic;
      \-adr12\        : in     std_logic;
      \-adr13\        : in     std_logic;
      \-adr14\        : in     std_logic;
      \-adr15\        : in     std_logic;
      \-adr16\        : in     std_logic;
      \-adr17\        : in     std_logic;
      \-adr18\        : in     std_logic;
      \-adr19\        : in     std_logic;
      \-adr1\         : in     std_logic;
      \-adr2\         : in     std_logic;
      \-adr3\         : in     std_logic;
      \-adr4\         : in     std_logic;
      \-adr5\         : in     std_logic;
      \-adr6\         : in     std_logic;
      \-adr7\         : in     std_logic;
      \-adr8\         : in     std_logic;
      \-adr9\         : in     std_logic;
      \-lmadr>ub\     : in     std_logic;
      \-lmadr>xbus\   : in     std_logic;
      uao1            : out    std_logic;
      uao10           : out    std_logic;
      uao11           : out    std_logic;
      uao12           : out    std_logic;
      uao13           : out    std_logic;
      uao14           : out    std_logic;
      uao15           : out    std_logic;
      uao16           : out    std_logic;
      uao17           : out    std_logic;
      uao2            : out    std_logic;
      uao3            : out    std_logic;
      uao4            : out    std_logic;
      uao5            : out    std_logic;
      uao6            : out    std_logic;
      uao7            : out    std_logic;
      uao8            : out    std_logic;
      uao9            : out    std_logic;
      xao0            : out    std_logic;
      xao1            : out    std_logic;
      xao10           : out    std_logic;
      xao11           : out    std_logic;
      xao12           : out    std_logic;
      xao13           : out    std_logic;
      xao14           : out    std_logic;
      xao15           : out    std_logic;
      xao16           : out    std_logic;
      xao17           : out    std_logic;
      xao18           : out    std_logic;
      xao19           : out    std_logic;
      xao2            : out    std_logic;
      xao3            : out    std_logic;
      xao4            : out    std_logic;
      xao5            : out    std_logic;
      xao6            : out    std_logic;
      xao7            : out    std_logic;
      xao8            : out    std_logic;
      xao9            : out    std_logic
    );
  end component;

  component cadr1_lmdata is
  port (
      \-lmbus enb\    : in     std_logic;
      \bus > lm\      : in     std_logic;
      bus0            : in     std_logic;
      bus1            : in     std_logic;
      bus10           : in     std_logic;
      bus11           : in     std_logic;
      bus12           : in     std_logic;
      bus13           : in     std_logic;
      bus14           : in     std_logic;
      bus15           : in     std_logic;
      bus16           : in     std_logic;
      bus17           : in     std_logic;
      bus18           : in     std_logic;
      bus19           : in     std_logic;
      bus2            : in     std_logic;
      bus20           : in     std_logic;
      bus21           : in     std_logic;
      bus22           : in     std_logic;
      bus23           : in     std_logic;
      bus24           : in     std_logic;
      bus25           : in     std_logic;
      bus26           : in     std_logic;
      bus27           : in     std_logic;
      bus28           : in     std_logic;
      bus29           : in     std_logic;
      bus3            : in     std_logic;
      bus30           : in     std_logic;
      bus31           : in     std_logic;
      bus4            : in     std_logic;
      bus5            : in     std_logic;
      bus6            : in     std_logic;
      bus7            : in     std_logic;
      bus8            : in     std_logic;
      bus9            : in     std_logic;
      mem10           : in     std_logic;
      mem11           : in     std_logic;
      mem18           : in     std_logic;
      mem19           : in     std_logic;
      mem20           : in     std_logic;
      mem21           : in     std_logic;
      mem22           : in     std_logic;
      mem23           : in     std_logic;
      mem30           : in     std_logic;
      mem31           : in     std_logic;
      mem6            : in     std_logic;
      mem7            : in     std_logic;
      mem8            : in     std_logic;
      mem9            : in     std_logic;
      mem0            : inout  std_logic;
      mem1            : inout  std_logic;
      mem12           : inout  std_logic;
      mem13           : inout  std_logic;
      mem14           : inout  std_logic;
      mem15           : inout  std_logic;
      mem16           : inout  std_logic;
      mem17           : inout  std_logic;
      mem2            : inout  std_logic;
      mem24           : inout  std_logic;
      mem25           : inout  std_logic;
      mem26           : inout  std_logic;
      mem27           : inout  std_logic;
      mem28           : inout  std_logic;
      mem29           : inout  std_logic;
      mem3            : inout  std_logic;
      mem4            : inout  std_logic;
      mem5            : inout  std_logic
    );
  end component;

  component cadr1_rbuf is
  port (
      \-bus>ub\       : in     std_logic;
      \-rbufwe\       : in     std_logic;
      \-ub read buffer\ : in     std_logic;
      \-ubpn0b\       : in     std_logic;
      \-ubpn1b\       : in     std_logic;
      \-ubpn2b\       : in     std_logic;
      \-ubpn3b\       : in     std_logic;
      bus0            : in     std_logic;
      bus1            : in     std_logic;
      bus10           : in     std_logic;
      bus11           : in     std_logic;
      bus12           : in     std_logic;
      bus13           : in     std_logic;
      bus14           : in     std_logic;
      bus15           : in     std_logic;
      bus16           : in     std_logic;
      bus17           : in     std_logic;
      bus18           : in     std_logic;
      bus19           : in     std_logic;
      bus2            : in     std_logic;
      bus20           : in     std_logic;
      bus21           : in     std_logic;
      bus22           : in     std_logic;
      bus23           : in     std_logic;
      bus24           : in     std_logic;
      bus25           : in     std_logic;
      bus26           : in     std_logic;
      bus27           : in     std_logic;
      bus28           : in     std_logic;
      bus29           : in     std_logic;
      bus3            : in     std_logic;
      bus30           : in     std_logic;
      bus31           : in     std_logic;
      bus4            : in     std_logic;
      bus5            : in     std_logic;
      bus6            : in     std_logic;
      bus7            : in     std_logic;
      bus8            : in     std_logic;
      bus9            : in     std_logic;
      rbuf16          : in     std_logic;
      rbuf17          : in     std_logic;
      rbuf18          : in     std_logic;
      rbuf19          : in     std_logic;
      rbuf20          : in     std_logic;
      rbuf21          : in     std_logic;
      rbuf22          : in     std_logic;
      rbuf23          : in     std_logic;
      rbuf24          : in     std_logic;
      rbuf25          : in     std_logic;
      rbuf26          : in     std_logic;
      rbuf27          : in     std_logic;
      rbuf28          : in     std_logic;
      rbuf29          : in     std_logic;
      rbuf30          : in     std_logic;
      rbuf31          : in     std_logic;
      udo0            : out    std_logic;
      udo1            : out    std_logic;
      udo10           : out    std_logic;
      udo11           : out    std_logic;
      udo12           : out    std_logic;
      udo13           : out    std_logic;
      udo14           : out    std_logic;
      udo15           : out    std_logic;
      udo2            : out    std_logic;
      udo3            : out    std_logic;
      udo4            : out    std_logic;
      udo5            : out    std_logic;
      udo6            : out    std_logic;
      udo7            : out    std_logic;
      udo8            : out    std_logic;
      udo9            : out    std_logic
    );
  end component;

  component cadr1_reqerr is
  port (
      \-adrpar\       : in     std_logic;
      \-db read status\ : in     std_logic;
      \-free\         : in     std_logic;
      \-int busy t80\ : in     std_logic;
      \-lmx grant\    : in     std_logic;
      \-nxm timeout\  : in     std_logic;
      \-reset err\    : in     std_logic;
      \-ub err drive\ : in     std_logic;
      \-ub invalid\   : in     std_logic;
      \-xao par even\ : in     std_logic;
      \bus par even\  : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \lm adr par error\ : in     std_logic;
      \lm par error\  : in     std_logic;
      \lmx grant a\   : in     std_logic;
      \mempar from lm\ : in     std_logic;
      \ub nxm error\  : in     std_logic;
      \ub xbus t100\  : in     std_logic;
      \unibus request\ : in     std_logic;
      \write through enb\ : in     std_logic;
      \xb nxm error\  : in     std_logic;
      \xb par error\  : in     std_logic;
      \xbus ignpar in\ : in     std_logic;
      \xbus par in\   : in     std_logic;
      \xbus request\  : in     std_logic;
      dbd0            : in     std_logic;
      dbd1            : in     std_logic;
      dbd2            : in     std_logic;
      dbd3            : in     std_logic;
      dbd4            : in     std_logic;
      dbd5            : in     std_logic;
      dbd6            : in     std_logic;
      dbd7            : in     std_logic;
      lmwr            : in     std_logic;
      xrd             : in     std_logic;
      \-xbus ignpar in\ : inout  std_logic;
      \ub map error\  : inout  std_logic;
      \-any par error\ : out    std_logic;
      \xbus par out\  : out    std_logic;
      udo0            : out    std_logic;
      udo1            : out    std_logic;
      udo2            : out    std_logic;
      udo3            : out    std_logic;
      udo4            : out    std_logic;
      udo5            : out    std_logic;
      udo6            : out    std_logic;
      udo7            : out    std_logic
    );
  end component;

  component cadr1_reqlm is
  port (
      \-adr17\        : in     std_logic;
      \-adr18\        : in     std_logic;
      \-adr19\        : in     std_logic;
      \-adr20\        : in     std_logic;
      \-adr21\        : in     std_logic;
      \-lm ub master\ : in     std_logic;
      \-lmub grant\   : in     std_logic;
      \-memrq\        : in     std_logic;
      \-ub to md\     : in     std_logic;
      \-ubx grant\    : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \int busy t100\ : in     std_logic;
      \int busy t80\  : in     std_logic;
      \lmub grant\    : in     std_logic;
      \lmx grant a\   : in     std_logic;
      \lmx grant\     : in     std_logic;
      \msyn in\       : in     std_logic;
      \nxm timeout\   : in     std_logic;
      \ssyn t150\     : in     std_logic;
      \ubx grant\     : in     std_logic;
      \unibus request\ : in     std_logic;
      \xbus ack in\   : in     std_logic;
      \xbus ignpar in\ : in     std_logic;
      lmrd            : in     std_logic;
      ubxrq           : in     std_logic;
      xrd             : in     std_logic;
      xwr             : in     std_logic;
      \-lmxrq\        : inout  std_logic;
      \-loadmd ack\   : inout  std_logic;
      \-xack\         : inout  std_logic;
      \adr=unibus\    : inout  std_logic;
      \ub md load\    : inout  std_logic;
      \xbus request\  : inout  std_logic;
      lmxrq           : inout  std_logic;
      xack            : inout  std_logic;
      \-lm grant\     : out    std_logic;
      \-lm ignpar\    : out    std_logic;
      \-lmack\        : out    std_logic;
      \-loadmd\       : out    std_logic;
      \-xbus request\ : out    std_logic;
      \lm memdrive enb\ : out    std_logic;
      \lmneedub (early)\ : out    std_logic;
      \loadmd ack\    : out    std_logic
    );
  end component;

  component cadr1_reqtim is
  port (
      \-debug timeout inh\ : in     std_logic;
      \int busy\      : in     std_logic;
      \select debug\  : in     std_logic;
      \timeout 0\     : in     std_logic;
      \timeout 1\     : in     std_logic;
      \timeout 2\     : in     std_logic;
      \timeout 3\     : in     std_logic;
      \vco cap2\      : in     std_logic;
      \hung timeout\  : inout  std_logic;
      \nxm timeout\   : inout  std_logic;
      \prom hung timeout\ : inout  std_logic;
      \prom nxm timeout\ : inout  std_logic;
      \prom unused\   : inout  std_logic;
      \vco cap1\      : inout  std_logic;
      \-hung timeout\ : out    std_logic;
      \-nxm timeout\  : out    std_logic;
      \unused timeout\ : out    std_logic
    );
  end component;

  component cadr1_requ is
  port (
      \-ub read xbus\ : in     std_logic;
      \-ub write xbus\ : in     std_logic;
      \-ubwr\         : in     std_logic;
      \-write through\ : in     std_logic;
      \debug ssyn\    : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \hi 15-30\      : in     std_logic;
      \intr ssyn\     : in     std_logic;
      \loadmd ack\    : in     std_logic;
      \msyn in\       : in     std_logic;
      \ub reg cyc t250\ : in     std_logic;
      \ub xbus t100\  : in     std_logic;
      \ubx grant a\   : in     std_logic;
      mapvalid        : in     std_logic;
      ubma17          : in     std_logic;
      ubma18          : in     std_logic;
      ubma19          : in     std_logic;
      ubma20          : in     std_logic;
      ubma21          : in     std_logic;
      ubwr            : in     std_logic;
      writeok         : in     std_logic;
      xack            : in     std_logic;
      \-uback\        : inout  std_logic;
      \-ubxrq\        : inout  std_logic;
      \ub xbus t0\    : inout  std_logic;
      ubxrq           : inout  std_logic;
      \-rbufwe\       : out    std_logic;
      \-ub invalid\   : out    std_logic;
      \-ub to md\     : out    std_logic;
      \ssyn out\      : out    std_logic
    );
  end component;

  component cadr1_requb is
  port (
      \-clk\          : in     std_logic;
      \db need ub\    : in     std_logic;
      \dbub master\   : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \int busy t100\ : in     std_logic;
      \lm ub master\  : in     std_logic;
      \lmneedub (early)\ : in     std_logic;
      \lmub grant\    : in     std_logic;
      \nxm timeout\   : in     std_logic;
      \ssyn in\       : in     std_logic;
      reset           : in     std_logic;
      \lm need ub\    : inout  std_logic;
      \ssyn t0\       : inout  std_logic;
      \ssyn t100\     : inout  std_logic;
      \unibus request\ : inout  std_logic;
      \-lm need ub\   : out    std_logic;
      \-unibus request\ : out    std_logic;
      \lmub rq\       : out    std_logic;
      \msyn out\      : out    std_logic;
      \ssyn t150\     : out    std_logic;
      \ssyn t200\     : out    std_logic;
      \ssyn t250\     : out    std_logic;
      \ssyn t50\      : out    std_logic
    );
  end component;

  component cadr1_rqsync is
  port (
      \-clk\          : in     std_logic;
      \-hung timeout\ : in     std_logic;
      \-lmxrq\        : in     std_logic;
      \-loadmd ack\   : in     std_logic;
      \-xbus request\ : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \hi 15-30\      : in     std_logic;
      \xbus busy in\  : in     std_logic;
      \xbus extrq in\ : in     std_logic;
      clk0            : in     std_logic;
      lmubrq          : in     std_logic;
      ubxrq           : in     std_logic;
      \-free\         : inout  std_logic;
      \-grant reset\  : inout  std_logic;
      \-lmub grant\   : inout  std_logic;
      \-lmubrqs\      : inout  std_logic;
      \-lmx grant\    : inout  std_logic;
      \-ubx grant\    : inout  std_logic;
      \-ubxrqs\       : inout  std_logic;
      \-xrqs\         : inout  std_logic;
      \int busy t40\  : inout  std_logic;
      \int busy t80\  : inout  std_logic;
      \int busy\      : inout  std_logic;
      \lmub grant set\ : inout  std_logic;
      \lmub grant\    : inout  std_logic;
      \lmx grant set\ : inout  std_logic;
      \ubx grant set\ : inout  std_logic;
      free            : inout  std_logic;
      lmubrqs         : inout  std_logic;
      ubxrqs          : inout  std_logic;
      xrqs            : inout  std_logic;
      \-int busy t80\ : out    std_logic;
      \grant reset\   : out    std_logic;
      \int busy t100\ : out    std_logic;
      \int busy t20\  : out    std_logic;
      \int busy t60\  : out    std_logic;
      \lmx grant a\   : out    std_logic;
      \lmx grant\     : out    std_logic;
      \ubx grant a\   : out    std_logic;
      \ubx grant\     : out    std_logic;
      \xbus extgrant out\ : out    std_logic
    );
  end component;

  component cadr1_uba is
  port (
      \-ub adr0\      : in     std_logic;
      \-ub adr10\     : in     std_logic;
      \-ub adr11\     : in     std_logic;
      \-ub adr12\     : in     std_logic;
      \-ub adr13\     : in     std_logic;
      \-ub adr14\     : in     std_logic;
      \-ub adr15\     : in     std_logic;
      \-ub adr16\     : in     std_logic;
      \-ub adr17\     : in     std_logic;
      \-ub adr1\      : in     std_logic;
      \-ub adr2\      : in     std_logic;
      \-ub adr3\      : in     std_logic;
      \-ub adr4\      : in     std_logic;
      \-ub adr5\      : in     std_logic;
      \-ub adr6\      : in     std_logic;
      \-ub adr7\      : in     std_logic;
      \-ub adr8\      : in     std_logic;
      \-ub adr9\      : in     std_logic;
      \-ub c1\        : in     std_logic;
      \-ubadrive\     : in     std_logic;
      \c1 in\         : in     std_logic;
      \c1 out\        : in     std_logic;
      uao1            : in     std_logic;
      uao10           : in     std_logic;
      uao11           : in     std_logic;
      uao12           : in     std_logic;
      uao13           : in     std_logic;
      uao14           : in     std_logic;
      uao15           : in     std_logic;
      uao16           : in     std_logic;
      uao17           : in     std_logic;
      uao2            : in     std_logic;
      uao3            : in     std_logic;
      uao4            : in     std_logic;
      uao5            : in     std_logic;
      uao6            : in     std_logic;
      uao7            : in     std_logic;
      uao8            : in     std_logic;
      uao9            : in     std_logic;
      uba0            : in     std_logic;
      uba1            : in     std_logic;
      uba10           : in     std_logic;
      uba11           : in     std_logic;
      uba12           : in     std_logic;
      uba13           : in     std_logic;
      uba14           : in     std_logic;
      uba15           : in     std_logic;
      uba16           : in     std_logic;
      uba17           : in     std_logic;
      uba2            : in     std_logic;
      uba3            : in     std_logic;
      uba4            : in     std_logic;
      uba5            : in     std_logic;
      uba6            : in     std_logic;
      uba7            : in     std_logic;
      uba8            : in     std_logic;
      uba9            : in     std_logic;
      \-uba 12\       : out    std_logic;
      \-uba 14\       : out    std_logic;
      \-uba 15\       : out    std_logic;
      \-uba 7\        : out    std_logic;
      \-uba 8\        : out    std_logic;
      \-uba 9\        : out    std_logic
    );
  end component;

  component cadr1_ubcyc is
  port (
      \-uba12\        : in     std_logic;
      \-uba14\        : in     std_logic;
      \-uba15\        : in     std_logic;
      \-uba7\         : in     std_logic;
      \-uba8\         : in     std_logic;
      \-uba9\         : in     std_logic;
      \-ubpn3a\       : in     std_logic;
      \c1 in\         : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \msyn in\       : in     std_logic;
      uba1            : in     std_logic;
      uba10           : in     std_logic;
      uba11           : in     std_logic;
      uba13           : in     std_logic;
      uba14           : in     std_logic;
      uba15           : in     std_logic;
      uba16           : in     std_logic;
      uba17           : in     std_logic;
      uba2            : in     std_logic;
      uba5            : in     std_logic;
      uba6            : in     std_logic;
      ubrd            : in     std_logic;
      ubwr            : in     std_logic;
      udi7            : in     std_logic;
      \-reset err\    : inout  std_logic;
      \-select interrupt\ : inout  std_logic;
      \-select page\  : inout  std_logic;
      \-select spy\   : inout  std_logic;
      \-ub read buffer\ : inout  std_logic;
      \-ub reg cyc t150\ : inout  std_logic;
      \-ub wr xbus\   : inout  std_logic;
      \-ub write buffer\ : inout  std_logic;
      \-write through enb\ : inout  std_logic;
      \-write through\ : inout  std_logic;
      \ub reg cyc t0\ : inout  std_logic;
      \ub reg cyc t150\ : inout  std_logic;
      \ub reg cyc t50\ : inout  std_logic;
      \ub reg write pulse\ : inout  std_logic;
      \ub17-14=map\   : inout  std_logic;
      \-intc drive\   : out    std_logic;
      \-load int ctl reg\ : out    std_logic;
      \-load int ctl2 reg\ : out    std_logic;
      \-select debug\ : out    std_logic;
      \-ub err drive\ : out    std_logic;
      \-ub read xbus\ : out    std_logic;
      \-ub write xbus\ : out    std_logic;
      \select page\   : out    std_logic;
      \ub reg cyc t100\ : out    std_logic;
      \ub reg cyc t200\ : out    std_logic;
      \ub reg cyc t250\ : out    std_logic;
      \write through enb\ : out    std_logic
    );
  end component;

  component cadr1_ubd is
  port (
      \-ubd0\         : in     std_logic;
      \-ubd10\        : in     std_logic;
      \-ubd11\        : in     std_logic;
      \-ubd12\        : in     std_logic;
      \-ubd13\        : in     std_logic;
      \-ubd14\        : in     std_logic;
      \-ubd15\        : in     std_logic;
      \-ubd1\         : in     std_logic;
      \-ubd2\         : in     std_logic;
      \-ubd3\         : in     std_logic;
      \-ubd4\         : in     std_logic;
      \-ubd5\         : in     std_logic;
      \-ubd6\         : in     std_logic;
      \-ubd7\         : in     std_logic;
      \-ubd8\         : in     std_logic;
      \-ubd9\         : in     std_logic;
      \-ubdrive\      : in     std_logic;
      \-udi > udo\    : in     std_logic;
      udi0            : in     std_logic;
      udi1            : in     std_logic;
      udi10           : in     std_logic;
      udi11           : in     std_logic;
      udi12           : in     std_logic;
      udi13           : in     std_logic;
      udi14           : in     std_logic;
      udi15           : in     std_logic;
      udi2            : in     std_logic;
      udi3            : in     std_logic;
      udi4            : in     std_logic;
      udi5            : in     std_logic;
      udi6            : in     std_logic;
      udi7            : in     std_logic;
      udi8            : in     std_logic;
      udi9            : in     std_logic;
      udo0            : inout  std_logic;
      udo1            : inout  std_logic;
      udo10           : inout  std_logic;
      udo11           : inout  std_logic;
      udo12           : inout  std_logic;
      udo13           : inout  std_logic;
      udo14           : inout  std_logic;
      udo15           : inout  std_logic;
      udo2            : inout  std_logic;
      udo3            : inout  std_logic;
      udo4            : inout  std_logic;
      udo5            : inout  std_logic;
      udo6            : inout  std_logic;
      udo7            : inout  std_logic;
      udo8            : inout  std_logic;
      udo9            : inout  std_logic
    );
  end component;

  component cadr1_ubintc is
  port (
      \-adr20\        : in     std_logic;
      \-adr21\        : in     std_logic;
      \-clk\          : in     std_logic;
      \-intc drive\   : in     std_logic;
      \-lmadr>xbus\   : in     std_logic;
      \-load int ctl reg\ : in     std_logic;
      \-load int ctl2 reg\ : in     std_logic;
      \-local enable\ : in     std_logic;
      \-reset\        : in     std_logic;
      \hi 15-30\      : in     std_logic;
      \local enable\  : in     std_logic;
      \unibus intr in\ : in     std_logic;
      \xbus intr in\  : in     std_logic;
      udi0            : in     std_logic;
      udi10           : in     std_logic;
      udi11           : in     std_logic;
      udi12           : in     std_logic;
      udi13           : in     std_logic;
      udi15           : in     std_logic;
      udi2            : in     std_logic;
      udi3            : in     std_logic;
      udi4            : in     std_logic;
      udi5            : in     std_logic;
      udi6            : in     std_logic;
      udi7            : in     std_logic;
      udi8            : in     std_logic;
      udi9            : in     std_logic;
      \-disable int grant\ : inout  std_logic;
      \-intr ssyn\    : inout  std_logic;
      \-ub int\       : inout  std_logic;
      \-xbus intr in\ : inout  std_logic;
      \enable ub ints\ : inout  std_logic;
      \int stops grants\ : inout  std_logic;
      \intr in\       : inout  std_logic;
      \intr ssyn\     : inout  std_logic;
      \ub int\        : inout  std_logic;
      \disable int grant\ : out    std_logic;
      \lm int\        : out    std_logic;
      level0          : out    std_logic;
      level1          : out    std_logic;
      udo0            : out    std_logic;
      udo1            : out    std_logic;
      udo10           : out    std_logic;
      udo11           : out    std_logic;
      udo12           : out    std_logic;
      udo13           : out    std_logic;
      udo14           : out    std_logic;
      udo15           : out    std_logic;
      udo2            : out    std_logic;
      udo3            : out    std_logic;
      udo4            : out    std_logic;
      udo5            : out    std_logic;
      udo6            : out    std_logic;
      udo7            : out    std_logic;
      udo8            : out    std_logic;
      udo9            : out    std_logic;
      xao20           : out    std_logic;
      xao21           : out    std_logic
    );
  end component;

  component cadr1_ubmap is
  port (
      \-ubmap > udo\  : in     std_logic;
      \-ubmapwe\      : in     std_logic;
      \select page\   : in     std_logic;
      mapvalid        : in     std_logic;
      uba1            : in     std_logic;
      uba10           : in     std_logic;
      uba11           : in     std_logic;
      uba12           : in     std_logic;
      uba13           : in     std_logic;
      uba2            : in     std_logic;
      uba3            : in     std_logic;
      uba4            : in     std_logic;
      ubma10          : in     std_logic;
      ubma11          : in     std_logic;
      ubma12          : in     std_logic;
      ubma13          : in     std_logic;
      ubma14          : in     std_logic;
      ubma15          : in     std_logic;
      ubma16          : in     std_logic;
      ubma17          : in     std_logic;
      ubma18          : in     std_logic;
      ubma19          : in     std_logic;
      ubma20          : in     std_logic;
      ubma21          : in     std_logic;
      ubma8           : in     std_logic;
      ubma9           : in     std_logic;
      udi0            : in     std_logic;
      udi1            : in     std_logic;
      udi10           : in     std_logic;
      udi11           : in     std_logic;
      udi12           : in     std_logic;
      udi13           : in     std_logic;
      udi14           : in     std_logic;
      udi15           : in     std_logic;
      udi2            : in     std_logic;
      udi3            : in     std_logic;
      udi4            : in     std_logic;
      udi5            : in     std_logic;
      udi6            : in     std_logic;
      udi7            : in     std_logic;
      udi8            : in     std_logic;
      udi9            : in     std_logic;
      writeok         : in     std_logic;
      \-ubpn0a\       : inout  std_logic;
      \-ubpn1a\       : inout  std_logic;
      \-ubpn2a\       : inout  std_logic;
      \-ubpn3a\       : inout  std_logic;
      \-ubpn0b\       : out    std_logic;
      \-ubpn1b\       : out    std_logic;
      \-ubpn2b\       : out    std_logic;
      \-ubpn3b\       : out    std_logic;
      udo0            : out    std_logic;
      udo1            : out    std_logic;
      udo10           : out    std_logic;
      udo11           : out    std_logic;
      udo12           : out    std_logic;
      udo13           : out    std_logic;
      udo14           : out    std_logic;
      udo15           : out    std_logic;
      udo2            : out    std_logic;
      udo3            : out    std_logic;
      udo4            : out    std_logic;
      udo5            : out    std_logic;
      udo6            : out    std_logic;
      udo7            : out    std_logic;
      udo8            : out    std_logic;
      udo9            : out    std_logic
    );
  end component;

  component cadr1_ubmast is
  port (
      \-db need ub\   : in     std_logic;
      \-dbub granted\ : in     std_logic;
      \-debug reset\  : in     std_logic;
      \-lm need ub\   : in     std_logic;
      \-lmub granted\ : in     std_logic;
      \-local enable\ : in     std_logic;
      \-npg in\       : in     std_logic;
      \-ub bbsy\      : in     std_logic;
      \-ub msyn\      : in     std_logic;
      \-ub sack\      : in     std_logic;
      \-ub ssyn\      : in     std_logic;
      \bbsy in\       : in     std_logic;
      \db need ub\    : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \msyn in\       : in     std_logic;
      \msyn out\      : in     std_logic;
      \npg1 in t100\  : in     std_logic;
      \npg1 in\       : in     std_logic;
      \npg2 in t100\  : in     std_logic;
      \npg2 in\       : in     std_logic;
      \sack in\       : in     std_logic;
      \ssyn in\       : in     std_logic;
      \ssyn out\      : in     std_logic;
      lmneedub        : in     std_logic;
      \-db bus req\   : inout  std_logic;
      \-db reset\     : inout  std_logic;
      \-db ub master\ : inout  std_logic;
      \-db ub selected\ : inout  std_logic;
      \-db ub set master\ : inout  std_logic;
      \-lm bus req\   : inout  std_logic;
      \-lm reset\     : inout  std_logic;
      \-lm ub master\ : inout  std_logic;
      \-lm ub selected\ : inout  std_logic;
      \-lm ub set master\ : inout  std_logic;
      \-npg1 out\     : inout  std_logic;
      \bus ready\     : inout  std_logic;
      \db ub granted\ : inout  std_logic;
      \db ub selected\ : inout  std_logic;
      \lm ub granted\ : inout  std_logic;
      \lm ub selected\ : inout  std_logic;
      \npg in\        : inout  std_logic;
      \npg1 out\      : inout  std_logic;
      \npg2 out\      : inout  std_logic;
      \-db ub granted\ : out    std_logic;
      \-lm ub granted\ : out    std_logic;
      \-npg out\      : out    std_logic;
      \bus req\       : out    std_logic;
      \db ub master\  : out    std_logic;
      \lm ub master\  : out    std_logic
    );
  end component;

  component cadr1_ubxa is
  port (
      \-ubaddr>xbus\  : in     std_logic;
      uba2            : in     std_logic;
      uba3            : in     std_logic;
      uba4            : in     std_logic;
      uba5            : in     std_logic;
      uba6            : in     std_logic;
      uba7            : in     std_logic;
      uba8            : in     std_logic;
      uba9            : in     std_logic;
      ubma10          : in     std_logic;
      ubma11          : in     std_logic;
      ubma12          : in     std_logic;
      ubma13          : in     std_logic;
      ubma14          : in     std_logic;
      ubma15          : in     std_logic;
      ubma16          : in     std_logic;
      ubma17          : in     std_logic;
      ubma18          : in     std_logic;
      ubma19          : in     std_logic;
      ubma20          : in     std_logic;
      ubma21          : in     std_logic;
      ubma8           : in     std_logic;
      ubma9           : in     std_logic;
      xao0            : out    std_logic;
      xao1            : out    std_logic;
      xao10           : out    std_logic;
      xao11           : out    std_logic;
      xao12           : out    std_logic;
      xao13           : out    std_logic;
      xao14           : out    std_logic;
      xao15           : out    std_logic;
      xao16           : out    std_logic;
      xao17           : out    std_logic;
      xao18           : out    std_logic;
      xao19           : out    std_logic;
      xao2            : out    std_logic;
      xao20           : out    std_logic;
      xao21           : out    std_logic;
      xao3            : out    std_logic;
      xao4            : out    std_logic;
      xao5            : out    std_logic;
      xao6            : out    std_logic;
      xao7            : out    std_logic;
      xao8            : out    std_logic;
      xao9            : out    std_logic
    );
  end component;

  component cadr1_uprior is
  port (
      \-clk\          : in     std_logic;
      \-disable int grant\ : in     std_logic;
      \-local enable\ : in     std_logic;
      \-npg in\       : in     std_logic;
      \-npg out\      : in     std_logic;
      \-ub br4\       : in     std_logic;
      \-ub br5\       : in     std_logic;
      \-ub br6\       : in     std_logic;
      \-ub br7\       : in     std_logic;
      \-ub init\      : in     std_logic;
      \-ub intr\      : in     std_logic;
      \-ub npr\       : in     std_logic;
      \bus req\       : in     std_logic;
      \grant timeout\ : in     std_logic;
      \hi 1-14\       : in     std_logic;
      \local enable\  : in     std_logic;
      \sack in\       : in     std_logic;
      \unibus init in\ : in     std_logic;
      \unibus intr in\ : in     std_logic;
      br4             : in     std_logic;
      br5             : in     std_logic;
      br6             : in     std_logic;
      br7             : in     std_logic;
      level0          : in     std_logic;
      level1          : in     std_logic;
      npr             : in     std_logic;
      reset           : in     std_logic;
      \-bg4o\         : inout  std_logic;
      \-bg5o\         : inout  std_logic;
      \-bg6o\         : inout  std_logic;
      \-bg7o\         : inout  std_logic;
      \-clear grant\  : inout  std_logic;
      \-npgo\         : inout  std_logic;
      \any grant dlyd\ : inout  std_logic;
      \any grant\     : inout  std_logic;
      \ub npg in\     : inout  std_logic;
      \ub npg out\    : inout  std_logic;
      bg4p            : inout  std_logic;
      bg5p            : inout  std_logic;
      bg6p            : inout  std_logic;
      bg7p            : inout  std_logic;
      br4d            : inout  std_logic;
      br5d            : inout  std_logic;
      br6d            : inout  std_logic;
      br7d            : inout  std_logic;
      npgp            : inout  std_logic;
      nprd            : inout  std_logic;
      sackd           : inout  std_logic;
      \-any grant dlyd\ : out    std_logic;
      \any int grant\ : out    std_logic;
      \ub bg4 in\     : out    std_logic;
      \ub bg5 in\     : out    std_logic;
      \ub bg6 in\     : out    std_logic;
      \ub bg7 in\     : out    std_logic;
      bg4o            : out    std_logic;
      bg5o            : out    std_logic;
      bg6o            : out    std_logic;
      bg7o            : out    std_logic;
      npgo            : out    std_logic
    );
  end component;

  component cadr1_wbuf is
  port (
      \-ubpn0a\       : in     std_logic;
      \-ubpn0b\       : in     std_logic;
      \-ubpn1a\       : in     std_logic;
      \-ubpn1b\       : in     std_logic;
      \-ubpn2a\       : in     std_logic;
      \-ubpn2b\       : in     std_logic;
      \-ubpn3a\       : in     std_logic;
      \-ubpn3b\       : in     std_logic;
      \-wbufwe\       : in     std_logic;
      udi0            : in     std_logic;
      udi1            : in     std_logic;
      udi10           : in     std_logic;
      udi11           : in     std_logic;
      udi12           : in     std_logic;
      udi13           : in     std_logic;
      udi14           : in     std_logic;
      udi15           : in     std_logic;
      udi2            : in     std_logic;
      udi3            : in     std_logic;
      udi4            : in     std_logic;
      udi5            : in     std_logic;
      udi6            : in     std_logic;
      udi7            : in     std_logic;
      udi8            : in     std_logic;
      udi9            : in     std_logic;
      wbuf0           : in     std_logic;
      wbuf1           : in     std_logic;
      wbuf10          : in     std_logic;
      wbuf11          : in     std_logic;
      wbuf12          : in     std_logic;
      wbuf13          : in     std_logic;
      wbuf14          : in     std_logic;
      wbuf15          : in     std_logic;
      wbuf2           : in     std_logic;
      wbuf3           : in     std_logic;
      wbuf4           : in     std_logic;
      wbuf5           : in     std_logic;
      wbuf6           : in     std_logic;
      wbuf7           : in     std_logic;
      wbuf8           : in     std_logic;
      wbuf9           : in     std_logic
    );
  end component;

  component cadr1_xa is
  port (
      \-lm power reset\ : in     std_logic;
      \-xaddrdrive\   : in     std_logic;
      \xaddr par out\ : in     std_logic;
      \xbus extgrant out\ : in     std_logic;
      \xbus request\  : in     std_logic;
      clk0            : in     std_logic;
      reset           : in     std_logic;
      xao0            : in     std_logic;
      xao1            : in     std_logic;
      xao10           : in     std_logic;
      xao11           : in     std_logic;
      xao12           : in     std_logic;
      xao13           : in     std_logic;
      xao14           : in     std_logic;
      xao15           : in     std_logic;
      xao16           : in     std_logic;
      xao17           : in     std_logic;
      xao18           : in     std_logic;
      xao19           : in     std_logic;
      xao2            : in     std_logic;
      xao20           : in     std_logic;
      xao21           : in     std_logic;
      xao3            : in     std_logic;
      xao4            : in     std_logic;
      xao5            : in     std_logic;
      xao6            : in     std_logic;
      xao7            : in     std_logic;
      xao8            : in     std_logic;
      xao9            : in     std_logic;
      \-xaddr par\    : inout  std_logic;
      \-xaddr0\       : inout  std_logic;
      \-xaddr10\      : inout  std_logic;
      \-xaddr11\      : inout  std_logic;
      \-xaddr12\      : inout  std_logic;
      \-xaddr13\      : inout  std_logic;
      \-xaddr14\      : inout  std_logic;
      \-xaddr15\      : inout  std_logic;
      \-xaddr16\      : inout  std_logic;
      \-xaddr17\      : inout  std_logic;
      \-xaddr18\      : inout  std_logic;
      \-xaddr19\      : inout  std_logic;
      \-xaddr1\       : inout  std_logic;
      \-xaddr20\      : inout  std_logic;
      \-xaddr21\      : inout  std_logic;
      \-xaddr2\       : inout  std_logic;
      \-xaddr3\       : inout  std_logic;
      \-xaddr4\       : inout  std_logic;
      \-xaddr5\       : inout  std_logic;
      \-xaddr6\       : inout  std_logic;
      \-xaddr7\       : inout  std_logic;
      \-xaddr8\       : inout  std_logic;
      \-xaddr9\       : inout  std_logic;
      \-xbus ack\     : inout  std_logic;
      \-xbus busy\    : inout  std_logic;
      \-xbus extgrant out\ : inout  std_logic;
      \-xbus extrq\   : inout  std_logic;
      \-xbus init\    : inout  std_logic;
      \-xbus intr\    : inout  std_logic;
      \-xbus power reset\ : inout  std_logic;
      \-xbus rq\      : inout  std_logic;
      \-xbus sync\    : inout  std_logic;
      \lm power reset\ : inout  std_logic;
      \xbus ack in\   : out    std_logic;
      \xbus busy in\  : out    std_logic;
      \xbus extrq in\ : out    std_logic;
      \xbus intr in\  : out    std_logic
    );
  end component;

  component cadr1_xapar is
  port (
      xao0            : in     std_logic;
      xao1            : in     std_logic;
      xao10           : in     std_logic;
      xao11           : in     std_logic;
      xao12           : in     std_logic;
      xao13           : in     std_logic;
      xao14           : in     std_logic;
      xao15           : in     std_logic;
      xao16           : in     std_logic;
      xao17           : in     std_logic;
      xao18           : in     std_logic;
      xao19           : in     std_logic;
      xao2            : in     std_logic;
      xao20           : in     std_logic;
      xao21           : in     std_logic;
      xao3            : in     std_logic;
      xao4            : in     std_logic;
      xao5            : in     std_logic;
      xao6            : in     std_logic;
      xao7            : in     std_logic;
      xao8            : in     std_logic;
      xao9            : in     std_logic;
      \xao par even\  : out    std_logic;
      \xao par odd\   : out    std_logic
    );
  end component;

  component cadr1_xbd is
  port (
      \-xb>bus\       : in     std_logic;
      xdi0            : in     std_logic;
      xdi1            : in     std_logic;
      xdi10           : in     std_logic;
      xdi11           : in     std_logic;
      xdi12           : in     std_logic;
      xdi13           : in     std_logic;
      xdi14           : in     std_logic;
      xdi15           : in     std_logic;
      xdi16           : in     std_logic;
      xdi17           : in     std_logic;
      xdi18           : in     std_logic;
      xdi19           : in     std_logic;
      xdi2            : in     std_logic;
      xdi20           : in     std_logic;
      xdi21           : in     std_logic;
      xdi22           : in     std_logic;
      xdi23           : in     std_logic;
      xdi24           : in     std_logic;
      xdi25           : in     std_logic;
      xdi26           : in     std_logic;
      xdi27           : in     std_logic;
      xdi28           : in     std_logic;
      xdi29           : in     std_logic;
      xdi3            : in     std_logic;
      xdi30           : in     std_logic;
      xdi31           : in     std_logic;
      xdi4            : in     std_logic;
      xdi5            : in     std_logic;
      xdi6            : in     std_logic;
      xdi7            : in     std_logic;
      xdi8            : in     std_logic;
      xdi9            : in     std_logic;
      bus0            : out    std_logic;
      bus1            : out    std_logic;
      bus10           : out    std_logic;
      bus11           : out    std_logic;
      bus12           : out    std_logic;
      bus13           : out    std_logic;
      bus14           : out    std_logic;
      bus15           : out    std_logic;
      bus16           : out    std_logic;
      bus17           : out    std_logic;
      bus18           : out    std_logic;
      bus19           : out    std_logic;
      bus2            : out    std_logic;
      bus20           : out    std_logic;
      bus21           : out    std_logic;
      bus22           : out    std_logic;
      bus23           : out    std_logic;
      bus24           : out    std_logic;
      bus25           : out    std_logic;
      bus26           : out    std_logic;
      bus27           : out    std_logic;
      bus28           : out    std_logic;
      bus29           : out    std_logic;
      bus3            : out    std_logic;
      bus30           : out    std_logic;
      bus31           : out    std_logic;
      bus4            : out    std_logic;
      bus5            : out    std_logic;
      bus6            : out    std_logic;
      bus7            : out    std_logic;
      bus8            : out    std_logic;
      bus9            : out    std_logic
    );
  end component;

  component cadr1_xd is
  port (
      \-xdrive\       : in     std_logic;
      \hi 15-30\      : in     std_logic;
      \xbus par out\  : in     std_logic;
      bus0            : in     std_logic;
      bus1            : in     std_logic;
      bus10           : in     std_logic;
      bus11           : in     std_logic;
      bus12           : in     std_logic;
      bus13           : in     std_logic;
      bus14           : in     std_logic;
      bus15           : in     std_logic;
      bus16           : in     std_logic;
      bus17           : in     std_logic;
      bus18           : in     std_logic;
      bus19           : in     std_logic;
      bus2            : in     std_logic;
      bus20           : in     std_logic;
      bus21           : in     std_logic;
      bus22           : in     std_logic;
      bus23           : in     std_logic;
      bus24           : in     std_logic;
      bus25           : in     std_logic;
      bus26           : in     std_logic;
      bus27           : in     std_logic;
      bus28           : in     std_logic;
      bus29           : in     std_logic;
      bus3            : in     std_logic;
      bus30           : in     std_logic;
      bus31           : in     std_logic;
      bus4            : in     std_logic;
      bus5            : in     std_logic;
      bus6            : in     std_logic;
      bus7            : in     std_logic;
      bus8            : in     std_logic;
      bus9            : in     std_logic;
      \-xbus ignpar\  : inout  std_logic;
      \-xbus par\     : inout  std_logic;
      \-xbus wr\      : inout  std_logic;
      \-xbus0\        : inout  std_logic;
      \-xbus10\       : inout  std_logic;
      \-xbus11\       : inout  std_logic;
      \-xbus12\       : inout  std_logic;
      \-xbus13\       : inout  std_logic;
      \-xbus14\       : inout  std_logic;
      \-xbus15\       : inout  std_logic;
      \-xbus16\       : inout  std_logic;
      \-xbus17\       : inout  std_logic;
      \-xbus18\       : inout  std_logic;
      \-xbus19\       : inout  std_logic;
      \-xbus1\        : inout  std_logic;
      \-xbus20\       : inout  std_logic;
      \-xbus21\       : inout  std_logic;
      \-xbus22\       : inout  std_logic;
      \-xbus23\       : inout  std_logic;
      \-xbus24\       : inout  std_logic;
      \-xbus25\       : inout  std_logic;
      \-xbus26\       : inout  std_logic;
      \-xbus27\       : inout  std_logic;
      \-xbus28\       : inout  std_logic;
      \-xbus29\       : inout  std_logic;
      \-xbus2\        : inout  std_logic;
      \-xbus30\       : inout  std_logic;
      \-xbus31\       : inout  std_logic;
      \-xbus3\        : inout  std_logic;
      \-xbus4\        : inout  std_logic;
      \-xbus5\        : inout  std_logic;
      \-xbus6\        : inout  std_logic;
      \-xbus7\        : inout  std_logic;
      \-xbus8\        : inout  std_logic;
      \-xbus9\        : inout  std_logic;
      \xbus ignpar in\ : out    std_logic;
      \xbus par in\   : out    std_logic;
      xdi0            : out    std_logic;
      xdi1            : out    std_logic;
      xdi10           : out    std_logic;
      xdi11           : out    std_logic;
      xdi12           : out    std_logic;
      xdi13           : out    std_logic;
      xdi14           : out    std_logic;
      xdi15           : out    std_logic;
      xdi16           : out    std_logic;
      xdi17           : out    std_logic;
      xdi18           : out    std_logic;
      xdi19           : out    std_logic;
      xdi2            : out    std_logic;
      xdi20           : out    std_logic;
      xdi21           : out    std_logic;
      xdi22           : out    std_logic;
      xdi23           : out    std_logic;
      xdi24           : out    std_logic;
      xdi25           : out    std_logic;
      xdi26           : out    std_logic;
      xdi27           : out    std_logic;
      xdi28           : out    std_logic;
      xdi29           : out    std_logic;
      xdi3            : out    std_logic;
      xdi30           : out    std_logic;
      xdi31           : out    std_logic;
      xdi4            : out    std_logic;
      xdi5            : out    std_logic;
      xdi6            : out    std_logic;
      xdi7            : out    std_logic;
      xdi8            : out    std_logic;
      xdi9            : out    std_logic
    );
  end component;

end package;
