library ieee;
use ieee.std_logic_1164.all;

entity cadr_clockd is
  port (
    \-srcpdlidx\    : in     std_logic;
    \-srcpdlptr\    : in     std_logic;
    \-tse1\         : in     std_logic;
    \-tse2\         : in     std_logic;
    \-tse3\         : in     std_logic;
    \-tse4\         : in     std_logic;
    \-wp1\          : in     std_logic;
    \-wp2\          : in     std_logic;
    \-wp3\          : in     std_logic;
    \-wp4\          : in     std_logic;
    clk1            : in     std_logic;
    clk2            : in     std_logic;
    clk3            : in     std_logic;
    clk4            : in     std_logic;
    hi1             : in     std_logic;
    hi10            : in     std_logic;
    hi11            : in     std_logic;
    hi12            : in     std_logic;
    hi2             : in     std_logic;
    hi3             : in     std_logic;
    hi4             : in     std_logic;
    hi5             : in     std_logic;
    hi6             : in     std_logic;
    hi7             : in     std_logic;
    hi8             : in     std_logic;
    hi9             : in     std_logic;
    lcry3           : in     std_logic;
    mclk1           : in     std_logic;
    reset           : in     std_logic;
    \-clk1\         : out    std_logic;
    \-clk2a\        : out    std_logic;
    \-clk2c\        : out    std_logic;
    \-clk3a\        : out    std_logic;
    \-clk3d\        : out    std_logic;
    \-clk3g\        : out    std_logic;
    \-clk4a\        : out    std_logic;
    \-clk4d\        : out    std_logic;
    \-clk4e\        : out    std_logic;
    \-lcry3\        : out    std_logic;
    \-mclk1\        : out    std_logic;
    \-reset\        : out    std_logic;
    \-upperhighok\  : out    std_logic;
    clk1a           : out    std_logic;
    clk2a           : out    std_logic;
    clk2b           : out    std_logic;
    clk2c           : out    std_logic;
    clk3a           : out    std_logic;
    clk3b           : out    std_logic;
    clk3c           : out    std_logic;
    clk3d           : out    std_logic;
    clk3e           : out    std_logic;
    clk3f           : out    std_logic;
    clk4a           : out    std_logic;
    clk4b           : out    std_logic;
    clk4c           : out    std_logic;
    clk4d           : out    std_logic;
    clk4e           : out    std_logic;
    clk4f           : out    std_logic;
    mclk1a          : out    std_logic;
    srcpdlidx       : out    std_logic;
    srcpdlptr       : out    std_logic;
    tse1a           : out    std_logic;
    tse1b           : out    std_logic;
    tse2            : out    std_logic;
    tse3a           : out    std_logic;
    tse4a           : out    std_logic;
    tse4b           : out    std_logic;
    wp1a            : out    std_logic;
    wp1b            : out    std_logic;
    wp2             : out    std_logic;
    wp3a            : out    std_logic;
    wp4a            : out    std_logic;
    wp4b            : out    std_logic;
    wp4c            : out    std_logic
  );
end entity;
