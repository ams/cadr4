library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn74260_tb is
end;

architecture testbench of sn74260_tb is

  signal g1a, g2a, g3a, g4a, g5a : std_logic;
  signal g1b, g2b, g3b, g4b, g5b : std_logic;
  signal g1y_n, g2y_n            : std_logic;

begin

  uut : sn74260 port map(
    g1a   => g1a,
    g2a   => g2a,
    g3a   => g3a,
    g4a   => g4a,
    g5a   => g5a,
    g1y_n => g1y_n,

    g1b   => g1b,
    g2b   => g2b,
    g3b   => g3b,
    g4b   => g4b,
    g5b   => g5b,
    g2y_n => g2y_n
    );

  process

    type pt is record
      i0, i1, i2, i3, i4 : std_logic;
      q                  : std_logic;
    end record;
    type pa is array (natural range <>) of pt;

    constant p : pa :=
      (('0', '0', '0', '0', '0', '1'),
       ('0', '0', '0', '0', '1', '0'),
       ('0', '0', '0', '1', '0', '0'),
       ('0', '0', '0', '1', '1', '0'),
       ('0', '0', '1', '0', '0', '0'),
       ('0', '0', '1', '0', '1', '0'),
       ('0', '0', '1', '1', '0', '0'),
       ('0', '0', '1', '1', '1', '0'),
       ('0', '1', '0', '0', '0', '0'),
       ('0', '1', '0', '0', '1', '0'),
       ('0', '1', '0', '1', '0', '0'),
       ('0', '1', '0', '1', '1', '0'),
       ('0', '1', '1', '0', '0', '0'),
       ('0', '1', '1', '0', '1', '0'),
       ('0', '1', '1', '1', '0', '0'),
       ('0', '1', '1', '1', '1', '0'),
       ('1', '0', '0', '0', '0', '0'),
       ('1', '0', '0', '0', '1', '0'),
       ('1', '0', '0', '1', '0', '0'),
       ('1', '0', '0', '1', '1', '0'),
       ('1', '0', '1', '0', '0', '0'),
       ('1', '0', '1', '0', '1', '0'),
       ('1', '0', '1', '1', '0', '0'),
       ('1', '0', '1', '1', '1', '0'),
       ('1', '1', '0', '0', '0', '0'),
       ('1', '1', '0', '0', '1', '0'),
       ('1', '1', '0', '1', '0', '0'),
       ('1', '1', '0', '1', '1', '0'),
       ('1', '1', '1', '0', '0', '0'),
       ('1', '1', '1', '0', '1', '0'),
       ('1', '1', '1', '1', '0', '0'),
       ('1', '1', '1', '1', '1', '0')
       );

  begin
    for i in p'range loop
      g1a <= p(i).i0; g2a <= p(i).i1; g3a <= p(i).i2; g4a <= p(i).i3; g5a <= p(i).i4;
      g1b <= p(i).i0; g2b <= p(i).i1; g3b <= p(i).i2; g4b <= p(i).i3; g5b <= p(i).i4;

      wait for 1 ns;

      assert g1y_n = p(i).q;
      assert g2y_n = p(i).q;
    end loop;

    wait;
  end process;

end;
