library ieee;
use ieee.std_logic_1164.all;

-- Dec 14 17:07:30 1980

package icmem_book is

  component clock1 is
    port ();
  end component;

  component clock2 is
    port ();
  end component;

  component debug is
    port ();
  end component;

  component icaps is
    port ();
  end component;

  component ictl is
    port ();
  end component;

  component iwrpar is
    port ();
  end component;

  component mbcpin is
    port ();
  end component;

  component mcpins is
    port ();
  end component;

  component olord1 is
    port ();
  end component;

  component olord2 is
    port ();
  end component;

  component opcs is
    port ();
  end component;

  component pctl is
    port ();
  end component;

  component prom0 is
    port ();
  end component;

  component prom1 is
    port ();
  end component;

  component iram00 is
    port ();
  end component;

  component iram01 is
    port ();
  end component;

  component iram02 is
    port ();
  end component;

  component iram03 is
    port ();
  end component;

  component iram10 is
    port ();
  end component;

  component iram11 is
    port ();
  end component;

  component iram12 is
    port ();
  end component;

  component iram13 is
    port ();
  end component;

  component iram20 is
    port ();
  end component;

  component iram21 is
    port ();
  end component;

  component iram22 is
    port ();
  end component;

  component iram23 is
    port ();
  end component;

  component iram30 is
    port ();
  end component;

  component iram31 is
    port ();
  end component;

  component iram32 is
    port ();
  end component;

  component iram33 is
    port ();
  end component;

  component spy0 is
    port ();
  end component;

  component spy4 is
    port ();
  end component;

  component stat is
    port ();
  end component;

end package;

