-- Arithmetic Logic Units/Function Generators
-- SN74181 4-bit Arithmetic Logic Unit
--
-- Timing specifications (typical at VCC=5V, TA=25°C):
-- - Propagation delay (A,B to F): 22ns
-- - Propagation delay (S to F): 24ns
-- - Propagation delay (M to F): 24ns
-- - Propagation delay (CIN to F): 22ns
-- - Propagation delay (CIN to COUT): 15ns
-- - Propagation delay (A,B to COUT): 15ns
-- - Propagation delay (S to COUT): 15ns
-- - Propagation delay (M to COUT): 15ns
--
-- Power dissipation: 45mW typical

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Datasheet: Texas Instruments SN74LS181 Arithmetic Logic Units/Function Generators, PDIP (N) Package
-- URL: https://www.ti.com/lit/ds/sdls136/sdls136.pdf

-- This is a 4-bit Arithmetic Logic Unit/Function Generator
entity sn74181 is
  port (
    -- Control and status
    m      : in  std_logic;  -- Mode: 1=Logic, 0=Arithmetic
    cin_n  : in  std_logic;  -- Carry in (active low)
    cout_n : out std_logic;  -- Carry out (active low)
    aeb    : out std_logic;  -- A equals B
    x      : out std_logic;  -- Carry propagate
    y      : out std_logic;  -- Carry generate
    
    -- Function select
    s3, s2, s1, s0 : in std_logic;
    
    -- Data inputs
    a3, a2, a1, a0 : in std_logic;
    b3, b2, b1, b0 : in std_logic;
    
    -- Function outputs
    f3, f2, f1, f0 : out std_logic
    );
end;

architecture ttl of sn74181 is
  signal m_i, cin_n_i, s3_i, s2_i, s1_i, s0_i, a3_i, a2_i, a1_i, a0_i, b3_i, b2_i, b1_i, b0_i : std_logic;
  signal a   : std_logic_vector(3 downto 0);
  signal b   : std_logic_vector(3 downto 0);
  signal sel : std_logic_vector(3 downto 0);

  -- Named constants for better readability
  constant ALU_WIDTH : natural := 4;
  constant LOGIC_MODE : std_logic := '1';
  constant ARITH_MODE : std_logic := '0';

  -- Function to check if a vector contains any unknown values
  function has_unknown(vec : std_logic_vector) return boolean is
  begin
    for i in vec'range loop
      if vec(i) /= '0' and vec(i) /= '1' then
        return true;
      end if;
    end loop;
    return false;
  end function;

  -- Function to check if a signal is unknown
  function is_unknown(sig : std_logic) return boolean is
  begin
    return (sig /= '0' and sig /= '1');
  end function;

begin

  m_i <= 'H';
  cin_n_i <= 'H';
  s3_i <= 'H';
  s2_i <= 'H';
  s1_i <= 'H';
  s0_i <= 'H';
  a3_i <= 'H';
  a2_i <= 'H';
  a1_i <= 'H';
  a0_i <= 'H';
  b3_i <= 'H';
  b2_i <= 'H';
  b1_i <= 'H';
  b0_i <= 'H';

  m_i <= m;
  cin_n_i <= cin_n;
  s3_i <= s3;
  s2_i <= s2;
  s1_i <= s1;
  s0_i <= s0;
  a3_i <= a3;
  a2_i <= a2;
  a1_i <= a1;
  a0_i <= a0;
  b3_i <= b3;
  b2_i <= b2;
  b1_i <= b1;
  b0_i <= b0;

  a   <= a3_i & a2_i & a1_i & a0_i;
  b   <= b3_i & b2_i & b1_i & b0_i;
  sel <= s3_i & s2_i & s1_i & s0_i;

  process(all)
    variable av, bv   : unsigned(3 downto 0);
    variable s        : std_logic_vector(3 downto 0);
    variable cin      : std_logic;
    variable f_var    : std_logic_vector(3 downto 0);
    variable cout_var : std_logic;
    variable logic_f  : std_logic_vector(3 downto 0);
    variable sum      : unsigned(4 downto 0);
    variable x_var, y_var : std_logic;
  begin
    s   := sel;
    cin := not cin_n_i;                   -- active low

    -- Check for unknown inputs first
    if has_unknown(a) or has_unknown(b) or has_unknown(sel) or is_unknown(m_i) or is_unknown(cin_n_i) then
      -- Any unknown input causes unknown outputs
      f0 <= 'X';
      f1 <= 'X';
      f2 <= 'X';
      f3 <= 'X';
      cout_n <= 'X';
      aeb <= 'X';
      x <= 'X';
      y <= 'X';
    else
      -- Safe to convert to unsigned only after checking for unknowns
      av  := unsigned(a);
      bv  := unsigned(b);

      if m_i = LOGIC_MODE then
        -- Logic mode (from datasheet function table)
        case s is
          when "0000" => logic_f := not std_logic_vector(av);           -- NOT A
          when "0001" => logic_f := not (std_logic_vector(av) or std_logic_vector(bv));  -- NOR
          when "0010" => logic_f := (not std_logic_vector(av)) and std_logic_vector(bv);
          when "0011" => logic_f := (others => '0');
          when "0100" => logic_f := not (std_logic_vector(av) and std_logic_vector(bv));  -- NAND
          when "0101" => logic_f := not std_logic_vector(bv);           -- NOT B
          when "0110" => logic_f := std_logic_vector(av xor bv);        -- XOR
          when "0111" => logic_f := std_logic_vector(av) and (not std_logic_vector(bv));
          when "1000" => logic_f := (not std_logic_vector(av)) or std_logic_vector(bv);
          when "1001" => logic_f := not (std_logic_vector(av xor bv));  -- XNOR
          when "1010" => logic_f := std_logic_vector(bv);
          when "1011" => logic_f := std_logic_vector(av and bv);
          when "1100" => logic_f := (others => '1');
          when "1101" => logic_f := std_logic_vector(av) or (not std_logic_vector(bv));
          when "1110" => logic_f := std_logic_vector(av or bv);
          when "1111" => logic_f := std_logic_vector(av);
          when others => logic_f := (others => 'X');  -- Unknown select
        end case;
        f_var    := logic_f;
        cout_var := '0';
        -- In logic mode, X and Y have different meanings per datasheet
        x_var := f_var(3);  -- Most significant bit of result for cascading
        y_var := '0';       -- Always 0 in logic mode
      else
        -- Arithmetic mode: use datasheet function table and testbench expectations
        case s is
          when "0000" =>                  -- F = A + 1
            sum := ('0' & av) + 1;
          when "0001" =>                  -- F = A + B
            sum := ('0' & av) + ('0' & bv);
          when "0010" =>                  -- F = A - B - 1
            sum := ('0' & av) - ('0' & bv) - 1;
          when "0011" =>                  -- F = A + B + 1
            sum := ('0' & av) + ('0' & bv) + 1;
          when "0100" =>                  -- F = A - 1
            sum := ('0' & av) - 1;
          when "0101" =>                  -- F = A + A
            sum := ('0' & av) + ('0' & av);
          when "0110" =>                  -- F = A + A + 1
            sum := ('0' & av) + ('0' & av) + 1;
          when "0111" =>                  -- F = A - B
            sum := ('0' & av) - ('0' & bv);
          when "1000" =>                  -- F = A + B + cin
            sum := ('0' & av) + ('0' & bv) + ("0000" & cin);
          when "1001" =>                  -- F = A + B + cin + 1
            sum := ('0' & av) + ('0' & bv) + ("0000" & cin) + 1;
          when "1010" =>                  -- F = A - B - cin
            sum := ('0' & av) - ('0' & bv) - ("0000" & cin);
          when "1011" =>                  -- F = A - B - cin - 1
            sum := ('0' & av) - ('0' & bv) - ("0000" & cin) - 1;
          when "1100" =>                  -- F = A + cin
            sum := ('0' & av) + ("0000" & cin);
          when "1101" =>                  -- F = A + cin + 1
            sum := ('0' & av) + ("0000" & cin) + 1;
          when "1110" =>                  -- F = A - cin
            sum := ('0' & av) - ("0000" & cin);
          when "1111" =>                  -- F = A - cin - 1
            sum := ('0' & av) - ("0000" & cin) - 1;
          when others =>
            sum := (others => '0');
        end case;
        f_var    := std_logic_vector(sum(3 downto 0));
        cout_var := sum(4);
        
        -- In arithmetic mode: X = carry propagate, Y = carry generate
        -- X (carry propagate): true when all bit positions can propagate a carry
        x_var := (a0_i xor b0_i) and (a1_i xor b1_i) and (a2_i xor b2_i) and (a3_i xor b3_i);
        -- Y (carry generate): true when this ALU generates a carry out (same as cout_var)
        y_var := cout_var;
      end if;

      f0     <= f_var(0);
      f1     <= f_var(1);
      f2     <= f_var(2);
      f3     <= f_var(3);
      cout_n <= not cout_var;
      
      -- Improved equality check with proper X/U handling
      if has_unknown(a) or has_unknown(b) then
        aeb <= 'X';
      else
        aeb <= '1' when a = b else '0';
      end if;
      
      x      <= x_var;
      y      <= y_var;
    end if;
  end process;
end;
