library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_vmas is
  port (
    vmasela     : in  std_logic;
    lc22        : in  std_logic;
    ob20        : in  std_logic;
    \-vmas20\   : out std_logic;
    lc23        : in  std_logic;
    ob21        : in  std_logic;
    \-vmas21\   : out std_logic;
    \-vmas22\   : out std_logic;
    ob22        : in  std_logic;
    lc24        : in  std_logic;
    \-vmas23\   : out std_logic;
    ob23        : in  std_logic;
    lc25        : in  std_logic;
    gnd         : in  std_logic;
    ob28        : in  std_logic;
    \-vmas28\   : out std_logic;
    ob29        : in  std_logic;
    \-vmas29\   : out std_logic;
    \-vmas30\   : out std_logic;
    ob30        : in  std_logic;
    \-vmas31\   : out std_logic;
    ob31        : in  std_logic;
    vmaselb     : in  std_logic;
    lc14        : in  std_logic;
    ob12        : in  std_logic;
    \-vmas12\   : out std_logic;
    lc15        : in  std_logic;
    ob13        : in  std_logic;
    \-vmas13\   : out std_logic;
    \-vmas14\   : out std_logic;
    ob14        : in  std_logic;
    lc16        : in  std_logic;
    \-vmas15\   : out std_logic;
    ob15        : in  std_logic;
    lc17        : in  std_logic;
    lc18        : in  std_logic;
    ob16        : in  std_logic;
    \-vmas16\   : out std_logic;
    lc19        : in  std_logic;
    ob17        : in  std_logic;
    \-vmas17\   : out std_logic;
    \-vmas18\   : out std_logic;
    ob18        : in  std_logic;
    lc20        : in  std_logic;
    \-vmas19\   : out std_logic;
    ob19        : in  std_logic;
    lc21        : in  std_logic;
    \-memstart\ : in  std_logic;
    \-vma12\    : in  std_logic;
    \-md12\     : in  std_logic;
    mapi12      : out std_logic;
    \-vma13\    : in  std_logic;
    \-md13\     : in  std_logic;
    mapi13      : out std_logic;
    mapi14      : out std_logic;
    \-md14\     : in  std_logic;
    \-vma14\    : in  std_logic;
    mapi15      : out std_logic;
    \-md15\     : in  std_logic;
    \-vma15\    : in  std_logic;
    \-vma16\    : in  std_logic;
    \-md16\     : in  std_logic;
    mapi16      : out std_logic;
    \-vma17\    : in  std_logic;
    \-md17\     : in  std_logic;
    mapi17      : out std_logic;
    mapi18      : out std_logic;
    \-md18\     : in  std_logic;
    \-vma18\    : in  std_logic;
    mapi19      : out std_logic;
    \-md19\     : in  std_logic;
    \-vma19\    : in  std_logic;
    \-vma20\    : in  std_logic;
    \-md20\     : in  std_logic;
    mapi20      : out std_logic;
    \-vma21\    : in  std_logic;
    \-md21\     : in  std_logic;
    mapi21      : out std_logic;
    mapi22      : out std_logic;
    \-md22\     : in  std_logic;
    \-vma22\    : in  std_logic;
    mapi23      : out std_logic;
    \-md23\     : in  std_logic;
    \-vma23\    : in  std_logic;
    lc2         : in  std_logic;
    ob0         : in  std_logic;
    \-vmas0\    : out std_logic;
    lc3         : in  std_logic;
    ob1         : in  std_logic;
    \-vmas1\    : out std_logic;
    \-vmas2\    : out std_logic;
    ob2         : in  std_logic;
    lc4         : in  std_logic;
    \-vmas3\    : out std_logic;
    ob3         : in  std_logic;
    lc5         : in  std_logic;
    \-vma8\     : in  std_logic;
    \-md8\      : in  std_logic;
    mapi8       : out std_logic;
    \-vma9\     : in  std_logic;
    \-md9\      : in  std_logic;
    mapi9       : out std_logic;
    mapi10      : out std_logic;
    \-md10\     : in  std_logic;
    \-vma10\    : in  std_logic;
    mapi11      : out std_logic;
    \-md11\     : in  std_logic;
    \-vma11\    : in  std_logic;
    lc10        : in  std_logic;
    ob8         : in  std_logic;
    \-vmas8\    : out std_logic;
    lc11        : in  std_logic;
    ob9         : in  std_logic;
    \-vmas9\    : out std_logic;
    \-vmas10\   : out std_logic;
    ob10        : in  std_logic;
    lc12        : in  std_logic;
    \-vmas11\   : out std_logic;
    ob11        : in  std_logic;
    lc13        : in  std_logic;
    lc6         : in  std_logic;
    ob4         : in  std_logic;
    \-vmas4\    : out std_logic;
    lc7         : in  std_logic;
    ob5         : in  std_logic;
    \-vmas5\    : out std_logic;
    \-vmas6\    : out std_logic;
    ob6         : in  std_logic;
    lc8         : in  std_logic;
    \-vmas7\    : out std_logic;
    ob7         : in  std_logic;
    lc9         : in  std_logic;
    ob24        : in  std_logic;
    \-vmas24\   : out std_logic;
    ob25        : in  std_logic;
    \-vmas25\   : out std_logic;
    \-vmas26\   : out std_logic;
    ob26        : in  std_logic;
    \-vmas27\   : out std_logic;
    ob27        : in  std_logic);
end;

architecture ttl of cadr_vmas is
begin
  vmas_1a27 : sn74s258 port map(sel => vmasela, d0 => lc22, d1 => ob20, dy => \-vmas20\, c0 => lc23, c1 => ob21, cy => \-vmas21\, by => \-vmas22\, b1 => ob22, b0 => lc24, ay => \-vmas23\, a1 => ob23, a0 => lc25, enb_n => gnd);
  vmas_1a29 : sn74s258 port map(sel => vmasela, d0 => gnd, d1 => ob28, dy => \-vmas28\, c0 => gnd, c1 => ob29, cy => \-vmas29\, by => \-vmas30\, b1 => ob30, b0 => gnd, ay => \-vmas31\, a1 => ob31, a0 => gnd, enb_n => gnd);
  vmas_1b26 : sn74s258 port map(sel => vmaselb, d0 => lc14, d1 => ob12, dy => \-vmas12\, c0 => lc15, c1 => ob13, cy => \-vmas13\, by => \-vmas14\, b1 => ob14, b0 => lc16, ay => \-vmas15\, a1 => ob15, a0 => lc17, enb_n => gnd);
  vmas_1b29 : sn74s258 port map(sel => vmasela, d0 => lc18, d1 => ob16, dy => \-vmas16\, c0 => lc19, c1 => ob17, cy => \-vmas17\, by => \-vmas18\, b1 => ob18, b0 => lc20, ay => \-vmas19\, a1 => ob19, a0 => lc21, enb_n => gnd);
  vmas_1c16 : sn74s258 port map(sel => \-memstart\, d0 => \-vma12\, d1 => \-md12\, dy => mapi12, c0 => \-vma13\, c1 => \-md13\, cy => mapi13, by => mapi14, b1 => \-md14\, b0 => \-vma14\, ay => mapi15, a1 => \-md15\, a0 => \-vma15\, enb_n => gnd);
  vmas_1c18 : sn74s258 port map(sel => \-memstart\, d0 => \-vma16\, d1 => \-md16\, dy => mapi16, c0 => \-vma17\, c1 => \-md17\, cy => mapi17, by => mapi18, b1 => \-md18\, b0 => \-vma18\, ay => mapi19, a1 => \-md19\, a0 => \-vma19\, enb_n => gnd);
  vmas_1c20 : sn74s258 port map(sel => \-memstart\, d0 => \-vma20\, d1 => \-md20\, dy => mapi20, c0 => \-vma21\, c1 => \-md21\, cy => mapi21, by => mapi22, b1 => \-md22\, b0 => \-vma22\, ay => mapi23, a1 => \-md23\, a0 => \-vma23\, enb_n => gnd);
  vmas_1c28 : sn74s258 port map(sel => vmaselb, d0 => lc2, d1 => ob0, dy => \-vmas0\, c0 => lc3, c1 => ob1, cy => \-vmas1\, by => \-vmas2\, b1 => ob2, b0 => lc4, ay => \-vmas3\, a1 => ob3, a0 => lc5, enb_n => gnd);
  vmas_1d19 : sn74s258 port map(sel => \-memstart\, d0 => \-vma8\, d1 => \-md8\, dy => mapi8, c0 => \-vma9\, c1 => \-md9\, cy => mapi9, by => mapi10, b1 => \-md10\, b0 => \-vma10\, ay => mapi11, a1 => \-md11\, a0 => \-vma11\, enb_n => gnd);
  vmas_1d30 : sn74s258 port map(sel => vmaselb, d0 => lc10, d1 => ob8, dy => \-vmas8\, c0 => lc11, c1 => ob9, cy => \-vmas9\, by => \-vmas10\, b1 => ob10, b0 => lc12, ay => \-vmas11\, a1 => ob11, a0 => lc13, enb_n => gnd);
  vmas_2b01 : sn74s258 port map(sel => vmaselb, d0 => lc6, d1 => ob4, dy => \-vmas4\, c0 => lc7, c1 => ob5, cy => \-vmas5\, by => \-vmas6\, b1 => ob6, b0 => lc8, ay => \-vmas7\, a1 => ob7, a0 => lc9, enb_n => gnd);
  vmas_2b04 : sn74s258 port map(sel => vmasela, d0 => gnd, d1 => ob24, dy => \-vmas24\, c0 => gnd, c1 => ob25, cy => \-vmas25\, by => \-vmas26\, b1 => ob26, b0 => gnd, ay => \-vmas27\, a1 => ob27, a0 => gnd, enb_n => gnd);
end architecture;
