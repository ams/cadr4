library ieee;
use ieee.std_logic_1164.all;

entity cadr_platch is
  port (
    \-pdldrive\ : in  std_logic;
    m15         : out std_logic;
    pdl15       : in  std_logic;
    pdl14       : in  std_logic;
    m14         : out std_logic;
    m13         : out std_logic;
    pdl13       : in  std_logic;
    pdl12       : in  std_logic;
    m12         : out std_logic;
    clk4a       : in  std_logic;
    m11         : out std_logic;
    pdl11       : in  std_logic;
    pdl10       : in  std_logic;
    m10         : out std_logic;
    m9          : out std_logic;
    pdl9        : in  std_logic;
    pdl8        : in  std_logic;
    m8          : out std_logic;
    m7          : out std_logic;
    pdl7        : in  std_logic;
    pdl6        : in  std_logic;
    m6          : out std_logic;
    m5          : out std_logic;
    pdl5        : in  std_logic;
    pdl4        : in  std_logic;
    m4          : out std_logic;
    m3          : out std_logic;
    pdl3        : in  std_logic;
    pdl2        : in  std_logic;
    m2          : out std_logic;
    m1          : out std_logic;
    pdl1        : in  std_logic;
    pdl0        : in  std_logic;
    m0          : out std_logic;
    m31         : out std_logic;
    pdl31       : in  std_logic;
    pdl30       : in  std_logic;
    m30         : out std_logic;
    m29         : out std_logic;
    pdl29       : in  std_logic;
    pdl28       : in  std_logic;
    m28         : out std_logic;
    m27         : out std_logic;
    pdl27       : in  std_logic;
    pdl26       : in  std_logic;
    m26         : out std_logic;
    m25         : out std_logic;
    pdl25       : in  std_logic;
    pdl24       : in  std_logic;
    m24         : out std_logic;
    m23         : out std_logic;
    pdl23       : in  std_logic;
    pdl22       : in  std_logic;
    m22         : out std_logic;
    m21         : out std_logic;
    pdl21       : in  std_logic;
    pdl20       : in  std_logic;
    m20         : out std_logic;
    m19         : out std_logic;
    pdl19       : in  std_logic;
    pdl18       : in  std_logic;
    m18         : out std_logic;
    m17         : out std_logic;
    pdl17       : in  std_logic;
    pdl16       : in  std_logic;
    m16         : out std_logic;
    pdlparity   : in  std_logic;
    mparity     : out std_logic
    );
end;
