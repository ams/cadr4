library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_dram0 is
  port (
    wp2         : in  std_logic;
    dispwr      : in  std_logic;
    \-dwea\     : out std_logic;
    nc418       : in  std_logic;
    nc419       : out std_logic;
    \-dadr10a\  : out std_logic;
    dadr10a     : out std_logic;
    ir22b       : in  std_logic;
    \-dadr9a\   : out std_logic;
    ir21b       : in  std_logic;
    \-dadr8a\   : out std_logic;
    ir20b       : in  std_logic;
    \-dadr7a\   : out std_logic;
    ir19b       : out std_logic;
    ir12b       : out std_logic;
    vmo19       : in  std_logic;
    ir9b        : in  std_logic;
    r0          : in  std_logic;
    dmask0      : in  std_logic;
    \-dmapbenb\ : in  std_logic;
    \-dadr0a\   : out std_logic;
    vmo18       : in  std_logic;
    ir8b        : in  std_logic;
    hi6         : in  std_logic;
    gnd         : in  std_logic;
    ir12        : in  std_logic;
    ir13        : in  std_logic;
    ir18b       : out std_logic;
    ir14        : in  std_logic;
    ir17b       : out std_logic;
    ir15        : in  std_logic;
    ir16b       : out std_logic;
    ir16        : in  std_logic;
    ir15b       : out std_logic;
    ir17        : in  std_logic;
    ir14b       : out std_logic;
    ir18        : in  std_logic;
    ir13b       : out std_logic;
    ir19        : in  std_logic;
    \-dadr1a\   : out std_logic;
    \-dadr2a\   : out std_logic;
    \-dadr3a\   : out std_logic;
    \-dadr4a\   : out std_logic;
    dpc5        : out std_logic;
    \-dadr5a\   : out std_logic;
    \-dadr6a\   : out std_logic;
    aa5         : in  std_logic;
    dpc4        : out std_logic;
    aa4         : in  std_logic;
    r3          : in  std_logic;
    dmask6      : in  std_logic;
    r6          : in  std_logic;
    dmask3      : in  std_logic;
    dpc3        : out std_logic;
    aa3         : in  std_logic;
    dpc2        : out std_logic;
    aa2         : in  std_logic;
    r2          : in  std_logic;
    hi4         : in  std_logic;
    dmask5      : in  std_logic;
    r5          : in  std_logic;
    dmask2      : in  std_logic;
    dpc1        : out std_logic;
    aa1         : in  std_logic;
    dpc0        : out std_logic;
    aa0         : in  std_logic;
    r1          : in  std_logic;
    dmask4      : in  std_logic;
    r4          : in  std_logic;
    dmask1      : in  std_logic);
end;

architecture ttl of cadr4_dram0 is
begin
  dram0_2f03 : sn74s37 port map(g1a     => wp2, g1b => dispwr, g1y => \-dwea\, g2a => '0', g2b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  dram0_2f21 : sn74s04 port map(g1a     => nc418, g1q_n => nc419, g2a => \-dadr10a\, g2q_n => dadr10a, g3a => ir22b, g3q_n => \-dadr10a\, g4q_n => \-dadr9a\, g4a => ir21b, g5q_n => \-dadr8a\, g5a => ir20b, g6q_n => \-dadr7a\, g6a => ir19b);
  dram0_2f24 : sn74s64 port map(d4      => ir12b, b2 => vmo19, a2 => ir9b, c3 => r0, b3 => dmask0, a3 => \-dmapbenb\, \out\ => \-dadr0a\, a1 => vmo18, b1 => ir8b, c4 => hi6, b4 => hi6, a4 => hi6);
  dram0_2f25 : sn74s241 port map(aenb_n => gnd, ain0 => ir12, bout3 => ir19b, ain1 => ir13, bout2 => ir18b, ain2 => ir14, bout1 => ir17b, ain3 => ir15, bout0 => ir16b, bin0 => ir16, aout3 => ir15b, bin1 => ir17, aout2 => ir14b, bin2 => ir18, aout1 => ir13b, bin3 => ir19, aout0 => ir12b, benb => hi6);
  dram0_2f26 : am93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc5, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa5);
  dram0_2f27 : am93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc5, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa5);
  dram0_2f28 : am93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc4, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa4);
  dram0_2f29 : am93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc4, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa4);
  dram0_2f30 : sn74s51 port map(g1a     => r3, g2a => ir18b, g2b => hi6, g2c => dmask6, g2d => r6, g2y => \-dadr6a\, g1y => \-dadr3a\, g1c => ir15b, g1d => hi6, g1b => dmask3);
  dram0_3f01 : am93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc3, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa3);
  dram0_3f02 : am93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc3, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa3);
  dram0_3f03 : am93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc2, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa2);
  dram0_3f04 : am93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc2, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa2);
  dram0_3f05 : sn74s51 port map(g1a     => r2, g2a => ir17b, g2b => hi4, g2c => dmask5, g2d => r5, g2y => \-dadr5a\, g1y => \-dadr2a\, g1c => ir14b, g1d => hi4, g1b => dmask2);
  dram0_3f06 : am93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc1, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa1);
  dram0_3f07 : am93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc1, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa1);
  dram0_3f08 : am93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc0, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa0);
  dram0_3f09 : am93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1 => \-dadr1a\, a2 => \-dadr2a\, a3 => \-dadr3a\, a4 => \-dadr4a\, do => dpc0, a5 => \-dadr5a\, a6 => \-dadr6a\, a7 => \-dadr7a\, a8 => \-dadr8a\, a9 => \-dadr9a\, we_n => \-dwea\, di => aa0);
  dram0_3f10 : sn74s51 port map(g1a     => r1, g2a => ir16b, g2b => hi4, g2c => dmask4, g2d => r4, g2y => \-dadr4a\, g1y => \-dadr1a\, g1c => ir13b, g1d => hi4, g1b => dmask1);
end architecture;
