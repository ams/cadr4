library ieee;
use ieee.std_logic_1164.all;

entity cadr1_ubintc is
  port (
    \-adr20\        : in     std_logic;
    \-adr21\        : in     std_logic;
    \-clk\          : in     std_logic;
    \-disable int grant\ : in     std_logic;
    \-intc drive\   : in     std_logic;
    \-intr ssyn\    : in     std_logic;
    \-lmadr>xbus\   : in     std_logic;
    \-load int ctl reg\ : in     std_logic;
    \-load int ctl2 reg\ : in     std_logic;
    \-local enable\ : in     std_logic;
    \-reset\        : in     std_logic;
    \-ub int\       : in     std_logic;
    \disable int grant\ : in     std_logic;
    \hi 15-30\      : in     std_logic;
    \intr ssyn\     : in     std_logic;
    \local enable\  : in     std_logic;
    \ub int\        : in     std_logic;
    \unibus intr in\ : in     std_logic;
    \xbus intr in\  : in     std_logic;
    udi0            : in     std_logic;
    udi10           : in     std_logic;
    udi11           : in     std_logic;
    udi12           : in     std_logic;
    udi13           : in     std_logic;
    udi15           : in     std_logic;
    udi2            : in     std_logic;
    udi3            : in     std_logic;
    udi4            : in     std_logic;
    udi5            : in     std_logic;
    udi6            : in     std_logic;
    udi7            : in     std_logic;
    udi8            : in     std_logic;
    udi9            : in     std_logic;
    \-xbus intr in\ : inout  std_logic;
    \enable ub ints\ : inout  std_logic;
    \int stops grants\ : inout  std_logic;
    \intr in\       : inout  std_logic;
    \lm int\        : out    std_logic;
    level0          : out    std_logic;
    level1          : out    std_logic;
    udo0            : out    std_logic;
    udo1            : out    std_logic;
    udo10           : out    std_logic;
    udo11           : out    std_logic;
    udo12           : out    std_logic;
    udo13           : out    std_logic;
    udo14           : out    std_logic;
    udo15           : out    std_logic;
    udo2            : out    std_logic;
    udo3            : out    std_logic;
    udo4            : out    std_logic;
    udo5            : out    std_logic;
    udo6            : out    std_logic;
    udo7            : out    std_logic;
    udo8            : out    std_logic;
    udo9            : out    std_logic;
    xao20           : out    std_logic;
    xao21           : out    std_logic
  );
end entity cadr1_ubintc;
