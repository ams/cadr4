library ieee;
use ieee.std_logic_1164.all;

entity cadr1_xa is
  port (
    \-lm power reset\ : in     std_logic;
    \-xaddr par\    : in     std_logic;
    \-xaddr0\       : in     std_logic;
    \-xaddr10\      : in     std_logic;
    \-xaddr11\      : in     std_logic;
    \-xaddr12\      : in     std_logic;
    \-xaddr13\      : in     std_logic;
    \-xaddr14\      : in     std_logic;
    \-xaddr15\      : in     std_logic;
    \-xaddr16\      : in     std_logic;
    \-xaddr17\      : in     std_logic;
    \-xaddr18\      : in     std_logic;
    \-xaddr19\      : in     std_logic;
    \-xaddr1\       : in     std_logic;
    \-xaddr20\      : in     std_logic;
    \-xaddr21\      : in     std_logic;
    \-xaddr2\       : in     std_logic;
    \-xaddr3\       : in     std_logic;
    \-xaddr4\       : in     std_logic;
    \-xaddr5\       : in     std_logic;
    \-xaddr6\       : in     std_logic;
    \-xaddr7\       : in     std_logic;
    \-xaddr8\       : in     std_logic;
    \-xaddr9\       : in     std_logic;
    \-xaddrdrive\   : in     std_logic;
    \-xbus ack\     : in     std_logic;
    \-xbus busy\    : in     std_logic;
    \-xbus extgrant out\ : in     std_logic;
    \-xbus extrq\   : in     std_logic;
    \-xbus init\    : in     std_logic;
    \-xbus intr\    : in     std_logic;
    \-xbus power reset\ : in     std_logic;
    \-xbus rq\      : in     std_logic;
    \-xbus sync\    : in     std_logic;
    \xaddr par out\ : in     std_logic;
    \xbus ack in\   : in     std_logic;
    \xbus busy in\  : in     std_logic;
    \xbus extgrant out\ : in     std_logic;
    \xbus extrq in\ : in     std_logic;
    \xbus intr in\  : in     std_logic;
    \xbus request\  : in     std_logic;
    clk0            : in     std_logic;
    reset           : in     std_logic;
    xao0            : in     std_logic;
    xao1            : in     std_logic;
    xao10           : in     std_logic;
    xao11           : in     std_logic;
    xao12           : in     std_logic;
    xao13           : in     std_logic;
    xao14           : in     std_logic;
    xao15           : in     std_logic;
    xao16           : in     std_logic;
    xao17           : in     std_logic;
    xao18           : in     std_logic;
    xao19           : in     std_logic;
    xao2            : in     std_logic;
    xao20           : in     std_logic;
    xao21           : in     std_logic;
    xao3            : in     std_logic;
    xao4            : in     std_logic;
    xao5            : in     std_logic;
    xao6            : in     std_logic;
    xao7            : in     std_logic;
    xao8            : in     std_logic;
    xao9            : in     std_logic;
    \lm power reset\ : inout  std_logic
  );
end entity cadr1_xa;
