library ieee;
use ieee.std_logic_1164.all;

entity busint_xbd is
  port (
    \-xb>bus\       : in     std_logic;
    xdi0            : in     std_logic;
    xdi1            : in     std_logic;
    xdi10           : in     std_logic;
    xdi11           : in     std_logic;
    xdi12           : in     std_logic;
    xdi13           : in     std_logic;
    xdi14           : in     std_logic;
    xdi15           : in     std_logic;
    xdi16           : in     std_logic;
    xdi17           : in     std_logic;
    xdi18           : in     std_logic;
    xdi19           : in     std_logic;
    xdi2            : in     std_logic;
    xdi20           : in     std_logic;
    xdi21           : in     std_logic;
    xdi22           : in     std_logic;
    xdi23           : in     std_logic;
    xdi24           : in     std_logic;
    xdi25           : in     std_logic;
    xdi26           : in     std_logic;
    xdi27           : in     std_logic;
    xdi28           : in     std_logic;
    xdi29           : in     std_logic;
    xdi3            : in     std_logic;
    xdi30           : in     std_logic;
    xdi31           : in     std_logic;
    xdi4            : in     std_logic;
    xdi5            : in     std_logic;
    xdi6            : in     std_logic;
    xdi7            : in     std_logic;
    xdi8            : in     std_logic;
    xdi9            : in     std_logic;
    bus0            : out    std_logic;
    bus1            : out    std_logic;
    bus10           : out    std_logic;
    bus11           : out    std_logic;
    bus12           : out    std_logic;
    bus13           : out    std_logic;
    bus14           : out    std_logic;
    bus15           : out    std_logic;
    bus16           : out    std_logic;
    bus17           : out    std_logic;
    bus18           : out    std_logic;
    bus19           : out    std_logic;
    bus2            : out    std_logic;
    bus20           : out    std_logic;
    bus21           : out    std_logic;
    bus22           : out    std_logic;
    bus23           : out    std_logic;
    bus24           : out    std_logic;
    bus25           : out    std_logic;
    bus26           : out    std_logic;
    bus27           : out    std_logic;
    bus28           : out    std_logic;
    bus29           : out    std_logic;
    bus3            : out    std_logic;
    bus30           : out    std_logic;
    bus31           : out    std_logic;
    bus4            : out    std_logic;
    bus5            : out    std_logic;
    bus6            : out    std_logic;
    bus7            : out    std_logic;
    bus8            : out    std_logic;
    bus9            : out    std_logic
  );
end entity busint_xbd;
