library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_7408 is
  port (
    g1b : in  std_logic;
    g1a : in  std_logic;
    g1q : out std_logic;
    g2b : in  std_logic;
    g2a : in  std_logic;
    g2q : out std_logic;
    g3a : in  std_logic;
    g3b : in  std_logic;
    g3q : out std_logic;
    g4q : out std_logic;
    g4a : in  std_logic;
    g4b : in  std_logic
    );
end ic_7408;

architecture ttl of ic_7408 is
begin

end ttl;
