library ieee;
use ieee.std_logic_1164.all;

entity cadr_mskg4 is
  port (
    \a=m\   : out std_logic;
    msk24   : out std_logic;
    msk25   : out std_logic;
    msk26   : out std_logic;
    msk27   : out std_logic;
    msk28   : out std_logic;
    msk29   : out std_logic;
    msk30   : out std_logic;
    msk31   : out std_logic;
    mskl0   : in  std_logic;
    mskl1   : in  std_logic;
    mskl2   : in  std_logic;
    mskl3   : in  std_logic;
    mskl4   : in  std_logic;
    gnd     : in  std_logic;
    mskr0   : in  std_logic;
    mskr1   : in  std_logic;
    mskr2   : in  std_logic;
    mskr3   : in  std_logic;
    mskr4   : in  std_logic;
    msk8    : out std_logic;
    msk9    : out std_logic;
    msk10   : out std_logic;
    msk11   : out std_logic;
    msk12   : out std_logic;
    msk13   : out std_logic;
    msk14   : out std_logic;
    msk15   : out std_logic;
    ir31    : in  std_logic;
    \-ir31\ : out std_logic;
    ir13    : in  std_logic;
    \-ir13\ : out std_logic;
    \-ir12\ : out std_logic;
    ir12    : in  std_logic;
    msk16   : out std_logic;
    msk17   : out std_logic;
    msk18   : out std_logic;
    msk19   : out std_logic;
    msk20   : out std_logic;
    msk21   : out std_logic;
    msk22   : out std_logic;
    msk23   : out std_logic;
    aeqm    : out std_logic;
    msk0    : out std_logic;
    msk1    : out std_logic;
    msk2    : out std_logic;
    msk3    : out std_logic;
    msk4    : out std_logic;
    msk5    : out std_logic;
    msk6    : out std_logic;
    msk7    : out std_logic);
end;
