library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_mctl is
  port (
    clk4e      : in  std_logic;
    wadr4      : in  std_logic;
    ir30       : in  std_logic;
    \-madr4a\  : out std_logic;
    \-madr4b\  : out std_logic;
    gnd        : in  std_logic;
    wadr0      : in  std_logic;
    ir26       : in  std_logic;
    \-madr0b\  : out std_logic;
    wadr1      : in  std_logic;
    ir27       : in  std_logic;
    \-madr1b\  : out std_logic;
    \-madr2b\  : out std_logic;
    ir28       : in  std_logic;
    wadr2      : in  std_logic;
    \-madr3b\  : out std_logic;
    ir29       : in  std_logic;
    wadr3      : in  std_logic;
    mmem15     : out std_logic;
    mmem14     : out std_logic;
    mmem13     : out std_logic;
    mmem12     : out std_logic;
    mmem11     : out std_logic;
    mmem10     : out std_logic;
    mmem9      : out std_logic;
    mmem8      : out std_logic;
    mmem7      : out std_logic;
    mmem6      : out std_logic;
    mmem5      : out std_logic;
    mmem4      : out std_logic;
    mmem3      : out std_logic;
    mmem2      : out std_logic;
    mmem1      : out std_logic;
    mmem0      : out std_logic;
    mpass      : out std_logic;
    tse4a      : in  std_logic;
    srcm       : out std_logic;
    hi2        : in  std_logic;
    \-ir31\    : in  std_logic;
    \-mpass\   : out std_logic;
    mpassl     : out std_logic;
    \-mpassm\  : out std_logic;
    \-mpassl\  : out std_logic;
    destmd     : in  std_logic;
    \-madr0a\  : out std_logic;
    \-madr1a\  : out std_logic;
    \-madr2a\  : out std_logic;
    \-madr3a\  : out std_logic;
    mmemparity : out std_logic;
    mmem31     : out std_logic;
    mmem30     : out std_logic;
    mmem29     : out std_logic;
    mmem28     : out std_logic;
    mmem27     : out std_logic;
    mmem26     : out std_logic;
    mmem25     : out std_logic;
    mmem24     : out std_logic;
    mmem23     : out std_logic;
    mmem22     : out std_logic;
    mmem21     : out std_logic;
    mmem20     : out std_logic;
    mmem19     : out std_logic;
    mmem18     : out std_logic;
    mmem17     : out std_logic;
    mmem16     : out std_logic;
    wp4b       : in  std_logic;
    \-mwpa\    : out std_logic;
    \-mwpb\    : out std_logic);
end;

architecture ttl of cadr_mctl is
  signal nc334 : std_logic;
  signal nc335 : std_logic;
  signal nc336 : std_logic;
  signal nc337 : std_logic;
  signal nc338 : std_logic;
  signal nc339 : std_logic;
  signal nc340 : std_logic;
begin
  mctl_4a16 : sn74s258 port map(sel => clk4e, d0 => wadr4, d1 => ir30, dy => \-madr4a\, c0 => nc335, c1 => nc336, cy => nc337, by => nc338, b1 => nc339, b0 => nc340, ay => \-madr4b\, a1 => ir30, a0 => wadr4, enb_n => gnd);
  mctl_4a18 : sn74s258 port map(sel => clk4e, d0 => wadr0, d1 => ir26, dy => \-madr0b\, c0 => wadr1, c1 => ir27, cy => \-madr1b\, by => \-madr2b\, b1 => ir28, b0 => wadr2, ay => \-madr3b\, a1 => ir29, a0 => wadr3, enb_n => gnd);
  mctl_4a19 : res20 port map(r2     => nc334, r3 => mmem15, r4 => mmem14, r5 => mmem13, r6 => mmem12, r7 => mmem11, r8 => mmem10, r9 => mmem9, r11 => mmem8, r12 => mmem7, r13 => mmem6, r14 => mmem5, r15 => mmem4, r16 => mmem3, r17 => mmem2, r18 => mmem1, r19 => mmem0);
  mctl_4b11 : sn74s11 port map(g1a  => mpass, g1b => tse4a, g3y => srcm, g3a => hi2, g3b => \-ir31\, g3c => \-mpass\, g1y => mpassl, g1c => \-ir31\, g2a => '0', g2b => '0', g2c => '0');
  mctl_4b12 : sn74s04 port map(g1a  => mpass, g1q_n => \-mpass\, g2a => '0', g3a => '0', g4a => '0', g5a => '0', g6a => '0');
  mctl_4b14 : sn74s10 port map(g1a  => mpass, g1b => tse4a, g2a => tse4a, g2b => \-ir31\, g2c => \-mpass\, g2y_n => \-mpassm\, g1y_n => \-mpassl\, g1c => \-ir31\, g3a => '0', g3b => '0', g3c => '0');
  mctl_4b18 : dm93s46 port map(a0   => ir26, b0 => wadr0, a1 => ir27, b1 => wadr1, a2 => ir28, b2 => wadr2, enb => hi2, eq => mpass, a3 => ir29, b3 => wadr3, a4 => ir30, b4 => wadr4, a5 => hi2, b5 => destmd);
  mctl_4b19 : sn74s258 port map(sel => clk4e, d0 => wadr0, d1 => ir26, dy => \-madr0a\, c0 => wadr1, c1 => ir27, cy => \-madr1a\, by => \-madr2a\, b1 => ir28, b0 => wadr2, ay => \-madr3a\, a1 => ir29, a0 => wadr3, enb_n => gnd);
  mctl_4b20 : res20 port map(r2     => mmemparity, r3 => mmem31, r4 => mmem30, r5 => mmem29, r6 => mmem28, r7 => mmem27, r8 => mmem26, r9 => mmem25, r11 => mmem24, r12 => mmem23, r13 => mmem22, r14 => mmem21, r15 => mmem20, r16 => mmem19, r17 => mmem18, r18 => mmem17, r19 => mmem16);
  mctl_4b22 : sn74s37 port map(g1a  => destmd, g1b => wp4b, g1y => \-mwpa\, g2a => destmd, g2b => wp4b, g2y => \-mwpb\, g3a => '0', g3b => '0', g4a => '0', g4b => '0');
end architecture;
