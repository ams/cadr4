library ieee;
use ieee.std_logic_1164.all;

entity cadr_pdlptr is
  port (
    \-srcpdlpop\ : in  std_logic;
    clk3f        : in  std_logic;
    ob8          : in  std_logic;
    ob9          : in  std_logic;
    \-destpdlp\  : in  std_logic;
    \-pdlcry7\   : out std_logic;
    pdlptr9      : out std_logic;
    pdlptr8      : out std_logic;
    \-destpdlx\  : in  std_logic;
    pdlidx6      : out std_logic;
    ob6          : in  std_logic;
    ob7          : in  std_logic;
    pdlidx7      : out std_logic;
    pdlidx8      : out std_logic;
    pdlidx9      : out std_logic;
    ob4          : in  std_logic;
    ob5          : in  std_logic;
    \-pdlcry3\   : out std_logic;
    pdlptr7      : out std_logic;
    pdlptr6      : out std_logic;
    pdlptr5      : out std_logic;
    pdlptr4      : out std_logic;
    pdlidx0      : out std_logic;
    ob0          : in  std_logic;
    ob1          : in  std_logic;
    pdlidx1      : out std_logic;
    ob2          : in  std_logic;
    pdlidx2      : out std_logic;
    pdlidx3      : out std_logic;
    ob3          : in  std_logic;
    pdlidx4      : out std_logic;
    pdlidx5      : out std_logic;
    \-pdlcnt\    : in  std_logic;
    pdlptr3      : out std_logic;
    pdlptr2      : out std_logic;
    pdlptr1      : out std_logic;
    pdlptr0      : out std_logic;
    \-ppdrive\   : out std_logic;
    mf0          : out std_logic;
    mf1          : out std_logic;
    mf2          : out std_logic;
    mf3          : out std_logic;
    pidrive      : out std_logic;
    mf8          : out std_logic;
    mf9          : out std_logic;
    mf10         : out std_logic;
    mf11         : out std_logic;
    mf4          : out std_logic;
    mf5          : out std_logic;
    mf6          : out std_logic;
    mf7          : out std_logic;
    srcpdlidx    : in  std_logic;
    tse4b        : in  std_logic;
    srcpdlptr    : in  std_logic
    );
end;
