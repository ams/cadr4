library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_ior is
  port (
    i12   : in  std_logic;
    ob12  : in  std_logic;
    iob12 : out std_logic;
    i13   : in  std_logic;
    ob13  : in  std_logic;
    iob13 : out std_logic;
    iob14 : out std_logic;
    i14   : in  std_logic;
    ob14  : in  std_logic;
    iob15 : out std_logic;
    i15   : in  std_logic;
    ob15  : in  std_logic;
    i8    : in  std_logic;
    ob8   : in  std_logic;
    iob8  : out std_logic;
    i9    : in  std_logic;
    ob9   : in  std_logic;
    iob9  : out std_logic;
    iob10 : out std_logic;
    i10   : in  std_logic;
    ob10  : in  std_logic;
    iob11 : out std_logic;
    i11   : in  std_logic;
    ob11  : in  std_logic;
    i4    : in  std_logic;
    ob4   : in  std_logic;
    iob4  : out std_logic;
    i5    : in  std_logic;
    ob5   : in  std_logic;
    iob5  : out std_logic;
    iob6  : out std_logic;
    i6    : in  std_logic;
    ob6   : in  std_logic;
    iob7  : out std_logic;
    i7    : in  std_logic;
    ob7   : in  std_logic;
    i0    : in  std_logic;
    ob0   : in  std_logic;
    iob0  : out std_logic;
    i1    : in  std_logic;
    ob1   : in  std_logic;
    iob1  : out std_logic;
    iob2  : out std_logic;
    i2    : in  std_logic;
    ob2   : in  std_logic;
    iob3  : out std_logic;
    i3    : in  std_logic;
    ob3   : in  std_logic;
    i20   : in  std_logic;
    ob20  : in  std_logic;
    iob20 : out std_logic;
    i21   : in  std_logic;
    ob21  : in  std_logic;
    iob21 : out std_logic;
    iob22 : out std_logic;
    i22   : in  std_logic;
    ob22  : in  std_logic;
    iob23 : out std_logic;
    i23   : in  std_logic;
    ob23  : in  std_logic;
    i16   : in  std_logic;
    ob16  : in  std_logic;
    iob16 : out std_logic;
    i17   : in  std_logic;
    ob17  : in  std_logic;
    iob17 : out std_logic;
    iob18 : out std_logic;
    i18   : in  std_logic;
    ob18  : in  std_logic;
    iob19 : out std_logic;
    i19   : in  std_logic;
    ob19  : in  std_logic;
    i44   : in  std_logic;
    iob44 : out std_logic;
    i45   : in  std_logic;
    iob45 : out std_logic;
    iob46 : out std_logic;
    i46   : in  std_logic;
    iob47 : out std_logic;
    i47   : in  std_logic;
    i40   : in  std_logic;
    iob40 : out std_logic;
    i41   : in  std_logic;
    iob41 : out std_logic;
    iob42 : out std_logic;
    i42   : in  std_logic;
    iob43 : out std_logic;
    i43   : in  std_logic;
    i36   : in  std_logic;
    iob36 : out std_logic;
    i37   : in  std_logic;
    iob37 : out std_logic;
    iob38 : out std_logic;
    i38   : in  std_logic;
    iob39 : out std_logic;
    i39   : in  std_logic;
    i32   : in  std_logic;
    iob32 : out std_logic;
    i33   : in  std_logic;
    iob33 : out std_logic;
    iob34 : out std_logic;
    i34   : in  std_logic;
    iob35 : out std_logic;
    i35   : in  std_logic;
    i28   : in  std_logic;
    iob28 : out std_logic;
    i29   : in  std_logic;
    iob29 : out std_logic;
    iob30 : out std_logic;
    i30   : in  std_logic;
    iob31 : out std_logic;
    i31   : in  std_logic;
    i24   : in  std_logic;
    ob24  : in  std_logic;
    iob24 : out std_logic;
    i25   : in  std_logic;
    ob25  : in  std_logic;
    iob25 : out std_logic;
    iob26 : out std_logic;
    i26   : in  std_logic;
    iob27 : out std_logic;
    i27   : in  std_logic);
end;

architecture ttl of cadr4_ior is
begin
  ior_3c06 : sn74s32 port map(g1a => i12, g1b => ob12, g1y => iob12, g2a => i13, g2b => ob13, g2y => iob13, g3y => iob14, g3a => i14, g3b => ob14, g4y => iob15, g4a => i15, g4b => ob15);
  ior_3c07 : sn74s32 port map(g1a => i8, g1b => ob8, g1y => iob8, g2a => i9, g2b => ob9, g2y => iob9, g3y => iob10, g3a => i10, g3b => ob10, g4y => iob11, g4a => i11, g4b => ob11);
  ior_3c08 : sn74s32 port map(g1a => i4, g1b => ob4, g1y => iob4, g2a => i5, g2b => ob5, g2y => iob5, g3y => iob6, g3a => i6, g3b => ob6, g4y => iob7, g4a => i7, g4b => ob7);
  ior_3c09 : sn74s32 port map(g1a => i0, g1b => ob0, g1y => iob0, g2a => i1, g2b => ob1, g2y => iob1, g3y => iob2, g3a => i2, g3b => ob2, g4y => iob3, g4a => i3, g4b => ob3);
  ior_3c16 : sn74s32 port map(g1a => i20, g1b => ob20, g1y => iob20, g2a => i21, g2b => ob21, g2y => iob21, g3y => iob22, g3a => i22, g3b => ob22, g4y => iob23, g4a => i23, g4b => ob23);
  ior_3c18 : sn74s32 port map(g1a => i16, g1b => ob16, g1y => iob16, g2a => i17, g2b => ob17, g2y => iob17, g3y => iob18, g3a => i18, g3b => ob18, g4y => iob19, g4a => i19, g4b => ob19);
  ior_3d08 : sn74s32 port map(g1a => i44, g1b => ob18, g1y => iob44, g2a => i45, g2b => ob19, g2y => iob45, g3y => iob46, g3a => i46, g3b => ob20, g4y => iob47, g4a => i47, g4b => ob21);
  ior_3d09 : sn74s32 port map(g1a => i40, g1b => ob14, g1y => iob40, g2a => i41, g2b => ob15, g2y => iob41, g3y => iob42, g3a => i42, g3b => ob16, g4y => iob43, g4a => i43, g4b => ob17);
  ior_3d10 : sn74s32 port map(g1a => i36, g1b => ob10, g1y => iob36, g2a => i37, g2b => ob11, g2y => iob37, g3y => iob38, g3a => i38, g3b => ob12, g4y => iob39, g4a => i39, g4b => ob13);
  ior_3d13 : sn74s32 port map(g1a => i32, g1b => ob6, g1y => iob32, g2a => i33, g2b => ob7, g2y => iob33, g3y => iob34, g3a => i34, g3b => ob8, g4y => iob35, g4a => i35, g4b => ob9);
  ior_3d14 : sn74s32 port map(g1a => i28, g1b => ob2, g1y => iob28, g2a => i29, g2b => ob3, g2y => iob29, g3y => iob30, g3a => i30, g3b => ob4, g4y => iob31, g4a => i31, g4b => ob5);
  ior_3d15 : sn74s32 port map(g1a => i24, g1b => ob24, g1y => iob24, g2a => i25, g2b => ob25, g2y => iob25, g3y => iob26, g3a => i26, g3b => ob0, g4y => iob27, g4a => i27, g4b => ob1);
end architecture;
