library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity helper_bus_monitor is 
    port (
      -- IPC bus (incremented PC, PC+1) - 14 bits
      ipc0    : in std_logic;
      ipc1    : in std_logic;
      ipc2    : in std_logic;
      ipc3    : in std_logic;
      ipc4    : in std_logic;
      ipc5    : in std_logic;
      ipc6    : in std_logic;
      ipc7    : in std_logic;
      ipc8    : in std_logic;
      ipc9    : in std_logic;
      ipc10   : in std_logic;
      ipc11   : in std_logic;
      ipc12   : in std_logic;
      ipc13   : in std_logic;
      -- IR bus (Instruction register) - 49 bits
      ir0     : in std_logic;
      ir1     : in std_logic;
      ir2     : in std_logic;
      ir3     : in std_logic;
      ir4     : in std_logic;
      ir5     : in std_logic;
      ir6     : in std_logic;
      ir7     : in std_logic;
      ir8     : in std_logic;
      ir9     : in std_logic;
      ir10    : in std_logic;
      ir11    : in std_logic;
      ir12    : in std_logic;
      ir13    : in std_logic;
      ir14    : in std_logic;
      ir15    : in std_logic;
      ir16    : in std_logic;
      ir17    : in std_logic;
      ir18    : in std_logic;
      ir19    : in std_logic;
      ir20    : in std_logic;
      ir21    : in std_logic;
      ir22    : in std_logic;
      ir23    : in std_logic;
      ir24    : in std_logic;
      ir25    : in std_logic;
      ir26    : in std_logic;
      ir27    : in std_logic;
      ir28    : in std_logic;
      ir29    : in std_logic;
      ir30    : in std_logic;
      ir31    : in std_logic;
      ir32    : in std_logic;
      ir33    : in std_logic;
      ir34    : in std_logic;
      ir35    : in std_logic;
      ir36    : in std_logic;
      ir37    : in std_logic;
      ir38    : in std_logic;
      ir39    : in std_logic;
      ir40    : in std_logic;
      ir41    : in std_logic;
      ir42    : in std_logic;
      ir43    : in std_logic;
      ir44    : in std_logic;
      ir45    : in std_logic;
      ir46    : in std_logic;
      ir47    : in std_logic;
      ir48    : in std_logic;
      -- NPC bus (Next PC) - 14 bits
      npc0    : in std_logic;
      npc1    : in std_logic;
      npc2    : in std_logic;
      npc3    : in std_logic;
      npc4    : in std_logic;
      npc5    : in std_logic;
      npc6    : in std_logic;
      npc7    : in std_logic;
      npc8    : in std_logic;
      npc9    : in std_logic;
      npc10   : in std_logic;
      npc11   : in std_logic;
      npc12   : in std_logic;
      npc13   : in std_logic;
      -- PC bus (Program counter) - 14 bits
      pc0     : in std_logic;
      pc1     : in std_logic;
      pc2     : in std_logic;
      pc3     : in std_logic;
      pc4     : in std_logic;
      pc5     : in std_logic;
      pc6     : in std_logic;
      pc7     : in std_logic;
      pc8     : in std_logic;
      pc9     : in std_logic;
      pc10    : in std_logic;
      pc11    : in std_logic;
      pc12    : in std_logic;
      pc13    : in std_logic;
      -- A bus (Address bus) - 31 bits
      a0      : in std_logic;
      a1      : in std_logic;
      a2      : in std_logic;
      a3      : in std_logic;
      a4      : in std_logic;
      a5      : in std_logic;
      a6      : in std_logic;
      a7      : in std_logic;
      a8      : in std_logic;
      a9      : in std_logic;
      a10     : in std_logic;
      a11     : in std_logic;
      a12     : in std_logic;
      a13     : in std_logic;
      a14     : in std_logic;
      a15     : in std_logic;
      a16     : in std_logic;
      a17     : in std_logic;
      a18     : in std_logic;
      a19     : in std_logic;
      a20     : in std_logic;
      a21     : in std_logic;
      a22     : in std_logic;
      a23     : in std_logic;
      a24     : in std_logic;
      a25     : in std_logic;
      a26     : in std_logic;
      a27     : in std_logic;
      a28     : in std_logic;
      a29     : in std_logic;
      a30     : in std_logic;
      -- L bus (L register) - 32 bits
      l0      : in std_logic;
      l1      : in std_logic;
      l2      : in std_logic;
      l3      : in std_logic;
      l4      : in std_logic;
      l5      : in std_logic;
      l6      : in std_logic;
      l7      : in std_logic;
      l8      : in std_logic;
      l9      : in std_logic;
      l10     : in std_logic;
      l11     : in std_logic;
      l12     : in std_logic;
      l13     : in std_logic;
      l14     : in std_logic;
      l15     : in std_logic;
      l16     : in std_logic;
      l17     : in std_logic;
      l18     : in std_logic;
      l19     : in std_logic;
      l20     : in std_logic;
      l21     : in std_logic;
      l22     : in std_logic;
      l23     : in std_logic;
      l24     : in std_logic;
      l25     : in std_logic;
      l26     : in std_logic;
      l27     : in std_logic;
      l28     : in std_logic;
      l29     : in std_logic;
      l30     : in std_logic;
      l31     : in std_logic;
      -- M bus (M register) - 32 bits
      m0      : in std_logic;
      m1      : in std_logic;
      m2      : in std_logic;
      m3      : in std_logic;
      m4      : in std_logic;
      m5      : in std_logic;
      m6      : in std_logic;
      m7      : in std_logic;
      m8      : in std_logic;
      m9      : in std_logic;
      m10     : in std_logic;
      m11     : in std_logic;
      m12     : in std_logic;
      m13     : in std_logic;
      m14     : in std_logic;
      m15     : in std_logic;
      m16     : in std_logic;
      m17     : in std_logic;
      m18     : in std_logic;
      m19     : in std_logic;
      m20     : in std_logic;
      m21     : in std_logic;
      m22     : in std_logic;
      m23     : in std_logic;
      m24     : in std_logic;
      m25     : in std_logic;
      m26     : in std_logic;
      m27     : in std_logic;
      m28     : in std_logic;
      m29     : in std_logic;
      m30     : in std_logic;
      m31     : in std_logic;
      -- OB bus (Output bus) - 32 bits
      ob0     : in std_logic;
      ob1     : in std_logic;
      ob2     : in std_logic;
      ob3     : in std_logic;
      ob4     : in std_logic;
      ob5     : in std_logic;
      ob6     : in std_logic;
      ob7     : in std_logic;
      ob8     : in std_logic;
      ob9     : in std_logic;
      ob10    : in std_logic;
      ob11    : in std_logic;
      ob12    : in std_logic;
      ob13    : in std_logic;
      ob14    : in std_logic;
      ob15    : in std_logic;
      ob16    : in std_logic;
      ob17    : in std_logic;
      ob18    : in std_logic;
      ob19    : in std_logic;
      ob20    : in std_logic;
      ob21    : in std_logic;
      ob22    : in std_logic;
      ob23    : in std_logic;
      ob24    : in std_logic;
      ob25    : in std_logic;
      ob26    : in std_logic;
      ob27    : in std_logic;
      ob28    : in std_logic;
      ob29    : in std_logic;
      ob30    : in std_logic;
      ob31    : in std_logic;
      -- I bus (Instruction bus) - 49 bits
      i0      : in std_logic;
      i1      : in std_logic;
      i2      : in std_logic;
      i3      : in std_logic;
      i4      : in std_logic;
      i5      : in std_logic;
      i6      : in std_logic;
      i7      : in std_logic;
      i8      : in std_logic;
      i9      : in std_logic;
      i10     : in std_logic;
      i11     : in std_logic;
      i12     : in std_logic;
      i13     : in std_logic;
      i14     : in std_logic;
      i15     : in std_logic;
      i16     : in std_logic;
      i17     : in std_logic;
      i18     : in std_logic;
      i19     : in std_logic;
      i20     : in std_logic;
      i21     : in std_logic;
      i22     : in std_logic;
      i23     : in std_logic;
      i24     : in std_logic;
      i25     : in std_logic;
      i26     : in std_logic;
      i27     : in std_logic;
      i28     : in std_logic;
      i29     : in std_logic;
      i30     : in std_logic;
      i31     : in std_logic;
      i32     : in std_logic;
      i33     : in std_logic;
      i34     : in std_logic;
      i35     : in std_logic;
      i36     : in std_logic;
      i37     : in std_logic;
      i38     : in std_logic;
      i39     : in std_logic;
      i40     : in std_logic;
      i41     : in std_logic;
      i42     : in std_logic;
      i43     : in std_logic;
      i44     : in std_logic;
      i45     : in std_logic;
      i46     : in std_logic;
      i47     : in std_logic;
      i48     : in std_logic;
      -- SPY bus - 16 bits
      spy0    : in std_logic;
      spy1    : in std_logic;
      spy2    : in std_logic;
      spy3    : in std_logic;
      spy4    : in std_logic;
      spy5    : in std_logic;
      spy6    : in std_logic;
      spy7    : in std_logic;
      spy8    : in std_logic;
      spy9    : in std_logic;
      spy10   : in std_logic;
      spy11   : in std_logic;
      spy12   : in std_logic;
      spy13   : in std_logic;
      spy14   : in std_logic;
      spy15   : in std_logic;
      -- MEM bus (Memory bus) - 32 bits
      mem0    : in std_logic;
      mem1    : in std_logic;
      mem2    : in std_logic;
      mem3    : in std_logic;
      mem4    : in std_logic;
      mem5    : in std_logic;
      mem6    : in std_logic;
      mem7    : in std_logic;
      mem8    : in std_logic;
      mem9    : in std_logic;
      mem10   : in std_logic;
      mem11   : in std_logic;
      mem12   : in std_logic;
      mem13   : in std_logic;
      mem14   : in std_logic;
      mem15   : in std_logic;
      mem16   : in std_logic;
      mem17   : in std_logic;
      mem18   : in std_logic;
      mem19   : in std_logic;
      mem20   : in std_logic;
      mem21   : in std_logic;
      mem22   : in std_logic;
      mem23   : in std_logic;
      mem24   : in std_logic;
      mem25   : in std_logic;
      mem26   : in std_logic;
      mem27   : in std_logic;
      mem28   : in std_logic;
      mem29   : in std_logic;
      mem30   : in std_logic;
      mem31   : in std_logic;
      -- AMEM bus (A memory bus) - 32 bits
      amem0   : in std_logic;
      amem1   : in std_logic;
      amem2   : in std_logic;
      amem3   : in std_logic;
      amem4   : in std_logic;
      amem5   : in std_logic;
      amem6   : in std_logic;
      amem7   : in std_logic;
      amem8   : in std_logic;
      amem9   : in std_logic;
      amem10  : in std_logic;
      amem11  : in std_logic;
      amem12  : in std_logic;
      amem13  : in std_logic;
      amem14  : in std_logic;
      amem15  : in std_logic;
      amem16  : in std_logic;
      amem17  : in std_logic;
      amem18  : in std_logic;
      amem19  : in std_logic;
      amem20  : in std_logic;
      amem21  : in std_logic;
      amem22  : in std_logic;
      amem23  : in std_logic;
      amem24  : in std_logic;
      amem25  : in std_logic;
      amem26  : in std_logic;
      amem27  : in std_logic;
      amem28  : in std_logic;
      amem29  : in std_logic;
      amem30  : in std_logic;
      amem31  : in std_logic;
      -- VMA bus (Virtual memory address) - 32 bits
      \-vma0\ : in std_logic;
      \-vma1\ : in std_logic;
      \-vma2\ : in std_logic;
      \-vma3\ : in std_logic;
      \-vma4\ : in std_logic;
      \-vma5\ : in std_logic;
      \-vma6\ : in std_logic;
      \-vma7\ : in std_logic;
      \-vma8\ : in std_logic;
      \-vma9\ : in std_logic;
      \-vma10\: in std_logic;
      \-vma11\: in std_logic;
      \-vma12\: in std_logic;
      \-vma13\: in std_logic;
      \-vma14\: in std_logic;
      \-vma15\: in std_logic;
      \-vma16\: in std_logic;
      \-vma17\: in std_logic;
      \-vma18\: in std_logic;
      \-vma19\: in std_logic;
      \-vma20\: in std_logic;
      \-vma21\: in std_logic;
      \-vma22\: in std_logic;
      \-vma23\: in std_logic;
      \-vma24\: in std_logic;
      \-vma25\: in std_logic;
      \-vma26\: in std_logic;
      \-vma27\: in std_logic;
      \-vma28\: in std_logic;
      \-vma29\: in std_logic;
      \-vma30\: in std_logic;
      \-vma31\: in std_logic;
      -- MD bus (Memory data) - 32 bits
      \-md0\  : in std_logic;
      \-md1\  : in std_logic;
      \-md2\  : in std_logic;
      \-md3\  : in std_logic;
      \-md4\  : in std_logic;
      \-md5\  : in std_logic;
      \-md6\  : in std_logic;
      \-md7\  : in std_logic;
      \-md8\  : in std_logic;
      \-md9\  : in std_logic;
      \-md10\ : in std_logic;
      \-md11\ : in std_logic;
      \-md12\ : in std_logic;
      \-md13\ : in std_logic;
      \-md14\ : in std_logic;
      \-md15\ : in std_logic;
      \-md16\ : in std_logic;
      \-md17\ : in std_logic;
      \-md18\ : in std_logic;
      \-md19\ : in std_logic;
      \-md20\ : in std_logic;
      \-md21\ : in std_logic;
      \-md22\ : in std_logic;
      \-md23\ : in std_logic;
      \-md24\ : in std_logic;
      \-md25\ : in std_logic;
      \-md26\ : in std_logic;
      \-md27\ : in std_logic;
      \-md28\ : in std_logic;
      \-md29\ : in std_logic;
      \-md30\ : in std_logic;
      \-md31\ : in std_logic;
      -- ALU bus - 33 bits
      alu0    : in std_logic;
      alu1    : in std_logic;
      alu2    : in std_logic;
      alu3    : in std_logic;
      alu4    : in std_logic;
      alu5    : in std_logic;
      alu6    : in std_logic;
      alu7    : in std_logic;
      alu8    : in std_logic;
      alu9    : in std_logic;
      alu10   : in std_logic;
      alu11   : in std_logic;
      alu12   : in std_logic;
      alu13   : in std_logic;
      alu14   : in std_logic;
      alu15   : in std_logic;
      alu16   : in std_logic;
      alu17   : in std_logic;
      alu18   : in std_logic;
      alu19   : in std_logic;
      alu20   : in std_logic;
      alu21   : in std_logic;
      alu22   : in std_logic;
      alu23   : in std_logic;
      alu24   : in std_logic;
      alu25   : in std_logic;
      alu26   : in std_logic;
      alu27   : in std_logic;
      alu28   : in std_logic;
      alu29   : in std_logic;
      alu30   : in std_logic;
      alu31   : in std_logic;
      alu32   : in std_logic;
      -- Q bus - 32 bits
      q0      : in std_logic;
      q1      : in std_logic;
      q2      : in std_logic;
      q3      : in std_logic;
      q4      : in std_logic;
      q5      : in std_logic;
      q6      : in std_logic;
      q7      : in std_logic;
      q8      : in std_logic;
      q9      : in std_logic;
      q10     : in std_logic;
      q11     : in std_logic;
      q12     : in std_logic;
      q13     : in std_logic;
      q14     : in std_logic;
      q15     : in std_logic;
      q16     : in std_logic;
      q17     : in std_logic;
      q18     : in std_logic;
      q19     : in std_logic;
      q20     : in std_logic;
      q21     : in std_logic;
      q22     : in std_logic;
      q23     : in std_logic;
      q24     : in std_logic;
      q25     : in std_logic;
      q26     : in std_logic;
      q27     : in std_logic;
      q28     : in std_logic;
      q29     : in std_logic;
      q30     : in std_logic;
      q31     : in std_logic;
      -- R bus - 32 bits
      r0      : in std_logic;
      r1      : in std_logic;
      r2      : in std_logic;
      r3      : in std_logic;
      r4      : in std_logic;
      r5      : in std_logic;
      r6      : in std_logic;
      r7      : in std_logic;
      r8      : in std_logic;
      r9      : in std_logic;
      r10     : in std_logic;
      r11     : in std_logic;
      r12     : in std_logic;
      r13     : in std_logic;
      r14     : in std_logic;
      r15     : in std_logic;
      r16     : in std_logic;
      r17     : in std_logic;
      r18     : in std_logic;
      r19     : in std_logic;
      r20     : in std_logic;
      r21     : in std_logic;
      r22     : in std_logic;
      r23     : in std_logic;
      r24     : in std_logic;
      r25     : in std_logic;
      r26     : in std_logic;
      r27     : in std_logic;
      r28     : in std_logic;
      r29     : in std_logic;
      r30     : in std_logic;
      r31     : in std_logic;
      -- AA bus - 18 bits
      aa0     : in std_logic;
      aa1     : in std_logic;
      aa2     : in std_logic;
      aa3     : in std_logic;
      aa4     : in std_logic;
      aa5     : in std_logic;
      aa6     : in std_logic;
      aa7     : in std_logic;
      aa8     : in std_logic;
      aa9     : in std_logic;
      aa10    : in std_logic;
      aa11    : in std_logic;
      aa12    : in std_logic;
      aa13    : in std_logic;
      aa14    : in std_logic;
      aa15    : in std_logic;
      aa16    : in std_logic;
      aa17    : in std_logic;
      -- DC bus - 10 bits
      dc0     : in std_logic;
      dc1     : in std_logic;
      dc2     : in std_logic;
      dc3     : in std_logic;
      dc4     : in std_logic;
      dc5     : in std_logic;
      dc6     : in std_logic;
      dc7     : in std_logic;
      dc8     : in std_logic;
      dc9     : in std_logic;
      -- DPC bus - 14 bits
      dpc0    : in std_logic;
      dpc1    : in std_logic;
      dpc2    : in std_logic;
      dpc3    : in std_logic;
      dpc4    : in std_logic;
      dpc5    : in std_logic;
      dpc6    : in std_logic;
      dpc7    : in std_logic;
      dpc8    : in std_logic;
      dpc9    : in std_logic;
      dpc10   : in std_logic;
      dpc11   : in std_logic;
      dpc12   : in std_logic;
      dpc13   : in std_logic;
      -- IWR bus - 49 bits
      iwr0    : in std_logic;
      iwr1    : in std_logic;
      iwr2    : in std_logic;
      iwr3    : in std_logic;
      iwr4    : in std_logic;
      iwr5    : in std_logic;
      iwr6    : in std_logic;
      iwr7    : in std_logic;
      iwr8    : in std_logic;
      iwr9    : in std_logic;
      iwr10   : in std_logic;
      iwr11   : in std_logic;
      iwr12   : in std_logic;
      iwr13   : in std_logic;
      iwr14   : in std_logic;
      iwr15   : in std_logic;
      iwr16   : in std_logic;
      iwr17   : in std_logic;
      iwr18   : in std_logic;
      iwr19   : in std_logic;
      iwr20   : in std_logic;
      iwr21   : in std_logic;
      iwr22   : in std_logic;
      iwr23   : in std_logic;
      iwr24   : in std_logic;
      iwr25   : in std_logic;
      iwr26   : in std_logic;
      iwr27   : in std_logic;
      iwr28   : in std_logic;
      iwr29   : in std_logic;
      iwr30   : in std_logic;
      iwr31   : in std_logic;
      iwr32   : in std_logic;
      iwr33   : in std_logic;
      iwr34   : in std_logic;
      iwr35   : in std_logic;
      iwr36   : in std_logic;
      iwr37   : in std_logic;
      iwr38   : in std_logic;
      iwr39   : in std_logic;
      iwr40   : in std_logic;
      iwr41   : in std_logic;
      iwr42   : in std_logic;
      iwr43   : in std_logic;
      iwr44   : in std_logic;
      iwr45   : in std_logic;
      iwr46   : in std_logic;
      iwr47   : in std_logic;
      iwr48   : in std_logic;
      -- LC bus - 26 bits
      lc0     : in std_logic;
      lc1     : in std_logic;
      lc2     : in std_logic;
      lc3     : in std_logic;
      lc4     : in std_logic;
      lc5     : in std_logic;
      lc6     : in std_logic;
      lc7     : in std_logic;
      lc8     : in std_logic;
      lc9     : in std_logic;
      lc10    : in std_logic;
      lc11    : in std_logic;
      lc12    : in std_logic;
      lc13    : in std_logic;
      lc14    : in std_logic;
      lc15    : in std_logic;
      lc16    : in std_logic;
      lc17    : in std_logic;
      lc18    : in std_logic;
      lc19    : in std_logic;
      lc20    : in std_logic;
      lc21    : in std_logic;
      lc22    : in std_logic;
      lc23    : in std_logic;
      lc24    : in std_logic;
      lc25    : in std_logic;
      -- MAPI bus - 16 bits (mapi8-mapi23)
      mapi8   : in std_logic;
      mapi9   : in std_logic;
      mapi10  : in std_logic;
      mapi11  : in std_logic;
      mapi12  : in std_logic;
      mapi13  : in std_logic;
      mapi14  : in std_logic;
      mapi15  : in std_logic;
      mapi16  : in std_logic;
      mapi17  : in std_logic;
      mapi18  : in std_logic;
      mapi19  : in std_logic;
      mapi20  : in std_logic;
      mapi21  : in std_logic;
      mapi22  : in std_logic;
      mapi23  : in std_logic;
      -- MSK bus - 32 bits
      msk0    : in std_logic;
      msk1    : in std_logic;
      msk2    : in std_logic;
      msk3    : in std_logic;
      msk4    : in std_logic;
      msk5    : in std_logic;
      msk6    : in std_logic;
      msk7    : in std_logic;
      msk8    : in std_logic;
      msk9    : in std_logic;
      msk10   : in std_logic;
      msk11   : in std_logic;
      msk12   : in std_logic;
      msk13   : in std_logic;
      msk14   : in std_logic;
      msk15   : in std_logic;
      msk16   : in std_logic;
      msk17   : in std_logic;
      msk18   : in std_logic;
      msk19   : in std_logic;
      msk20   : in std_logic;
      msk21   : in std_logic;
      msk22   : in std_logic;
      msk23   : in std_logic;
      msk24   : in std_logic;
      msk25   : in std_logic;
      msk26   : in std_logic;
      msk27   : in std_logic;
      msk28   : in std_logic;
      msk29   : in std_logic;
      msk30   : in std_logic;
      msk31   : in std_logic;
      -- OPC bus - 14 bits
      opc0    : in std_logic;
      opc1    : in std_logic;
      opc2    : in std_logic;
      opc3    : in std_logic;
      opc4    : in std_logic;
      opc5    : in std_logic;
      opc6    : in std_logic;
      opc7    : in std_logic;
      opc8    : in std_logic;
      opc9    : in std_logic;
      opc10   : in std_logic;
      opc11   : in std_logic;
      opc12   : in std_logic;
      opc13   : in std_logic;
      -- SPC bus - 19 bits
      spc0    : in std_logic;
      spc1    : in std_logic;
      spc2    : in std_logic;
      spc3    : in std_logic;
      spc4    : in std_logic;
      spc5    : in std_logic;
      spc6    : in std_logic;
      spc7    : in std_logic;
      spc8    : in std_logic;
      spc9    : in std_logic;
      spc10   : in std_logic;
      spc11   : in std_logic;
      spc12   : in std_logic;
      spc13   : in std_logic;
      spc14   : in std_logic;
      spc15   : in std_logic;
      spc16   : in std_logic;
      spc17   : in std_logic;
      spc18   : in std_logic;
      -- WADR bus - 10 bits
      wadr0   : in std_logic;
      wadr1   : in std_logic;
      wadr2   : in std_logic;
      wadr3   : in std_logic;
      wadr4   : in std_logic;
      wadr5   : in std_logic;
      wadr6   : in std_logic;
      wadr7   : in std_logic;
      wadr8   : in std_logic;
      wadr9   : in std_logic
    );
  end entity;

  architecture structural of helper_bus_monitor is
    signal ipc : std_logic_vector(13 downto 0);
    signal ir : std_logic_vector(48 downto 0);
    signal npc : std_logic_vector(13 downto 0);
    signal pc : std_logic_vector(13 downto 0);
    signal a : std_logic_vector(30 downto 0);
    signal l : std_logic_vector(31 downto 0);
    signal m : std_logic_vector(31 downto 0);
    signal ob : std_logic_vector(31 downto 0);
    signal i : std_logic_vector(48 downto 0);
    signal spy : std_logic_vector(15 downto 0);
    signal mem : std_logic_vector(31 downto 0);
    signal amem : std_logic_vector(31 downto 0);
    signal vma : std_logic_vector(31 downto 0);
    signal md : std_logic_vector(31 downto 0);
    signal \-vma\ : std_logic_vector(31 downto 0);
    signal \-md\ : std_logic_vector(31 downto 0);
    signal alu : std_logic_vector(32 downto 0);
    signal q : std_logic_vector(31 downto 0);
    signal r : std_logic_vector(31 downto 0);
    signal aa : std_logic_vector(17 downto 0);
    signal dc : std_logic_vector(9 downto 0);
    signal dpc : std_logic_vector(13 downto 0);
    signal iwr : std_logic_vector(48 downto 0);
    signal lc : std_logic_vector(25 downto 0);
    signal mapi : std_logic_vector(15 downto 0);
    signal msk : std_logic_vector(31 downto 0);
    signal opc : std_logic_vector(13 downto 0);
    signal spc : std_logic_vector(18 downto 0);
    signal wadr : std_logic_vector(9 downto 0);
  begin
    ipc <= ipc13 & ipc12 & ipc11 & ipc10 & ipc9 & ipc8 & ipc7 & ipc6 & ipc5 & ipc4 & ipc3 & ipc2 & ipc1 & ipc0;
    ir <= ir48 & ir47 & ir46 & ir45 & ir44 & ir43 & ir42 & ir41 & ir40 & ir39 & ir38 & ir37 & ir36 & ir35 & ir34 & ir33 & ir32 & ir31 & ir30 & ir29 & ir28 & ir27 & ir26 & ir25 & ir24 & ir23 & ir22 & ir21 & ir20 & ir19 & ir18 & ir17 & ir16 & ir15 & ir14 & ir13 & ir12 & ir11 & ir10 & ir9 & ir8 & ir7 & ir6 & ir5 & ir4 & ir3 & ir2 & ir1 & ir0;
    npc <= npc13 & npc12 & npc11 & npc10 & npc9 & npc8 & npc7 & npc6 & npc5 & npc4 & npc3 & npc2 & npc1 & npc0;
    pc <= pc13 & pc12 & pc11 & pc10 & pc9 & pc8 & pc7 & pc6 & pc5 & pc4 & pc3 & pc2 & pc1 & pc0;
    a <= a30 & a29 & a28 & a27 & a26 & a25 & a24 & a23 & a22 & a21 & a20 & a19 & a18 & a17 & a16 & a15 & a14 & a13 & a12 & a11 & a10 & a9 & a8 & a7 & a6 & a5 & a4 & a3 & a2 & a1 & a0;
    l <= l31 & l30 & l29 & l28 & l27 & l26 & l25 & l24 & l23 & l22 & l21 & l20 & l19 & l18 & l17 & l16 & l15 & l14 & l13 & l12 & l11 & l10 & l9 & l8 & l7 & l6 & l5 & l4 & l3 & l2 & l1 & l0;
    m <= m31 & m30 & m29 & m28 & m27 & m26 & m25 & m24 & m23 & m22 & m21 & m20 & m19 & m18 & m17 & m16 & m15 & m14 & m13 & m12 & m11 & m10 & m9 & m8 & m7 & m6 & m5 & m4 & m3 & m2 & m1 & m0;
    ob <= ob31 & ob30 & ob29 & ob28 & ob27 & ob26 & ob25 & ob24 & ob23 & ob22 & ob21 & ob20 & ob19 & ob18 & ob17 & ob16 & ob15 & ob14 & ob13 & ob12 & ob11 & ob10 & ob9 & ob8 & ob7 & ob6 & ob5 & ob4 & ob3 & ob2 & ob1 & ob0;
    i <= i48 & i47 & i46 & i45 & i44 & i43 & i42 & i41 & i40 & i39 & i38 & i37 & i36 & i35 & i34 & i33 & i32 & i31 & i30 & i29 & i28 & i27 & i26 & i25 & i24 & i23 & i22 & i21 & i20 & i19 & i18 & i17 & i16 & i15 & i14 & i13 & i12 & i11 & i10 & i9 & i8 & i7 & i6 & i5 & i4 & i3 & i2 & i1 & i0;
    spy <= spy15 & spy14 & spy13 & spy12 & spy11 & spy10 & spy9 & spy8 & spy7 & spy6 & spy5 & spy4 & spy3 & spy2 & spy1 & spy0;
    mem <= mem31 & mem30 & mem29 & mem28 & mem27 & mem26 & mem25 & mem24 & mem23 & mem22 & mem21 & mem20 & mem19 & mem18 & mem17 & mem16 & mem15 & mem14 & mem13 & mem12 & mem11 & mem10 & mem9 & mem8 & mem7 & mem6 & mem5 & mem4 & mem3 & mem2 & mem1 & mem0;
    amem <= amem31 & amem30 & amem29 & amem28 & amem27 & amem26 & amem25 & amem24 & amem23 & amem22 & amem21 & amem20 & amem19 & amem18 & amem17 & amem16 & amem15 & amem14 & amem13 & amem12 & amem11 & amem10 & amem9 & amem8 & amem7 & amem6 & amem5 & amem4 & amem3 & amem2 & amem1 & amem0;
    \-vma\ <= \-vma31\ & \-vma30\ & \-vma29\ & \-vma28\ & \-vma27\ & \-vma26\ & \-vma25\ & \-vma24\ & \-vma23\ & \-vma22\ & \-vma21\ & \-vma20\ & \-vma19\ & \-vma18\ & \-vma17\ & \-vma16\ & \-vma15\ & \-vma14\ & \-vma13\ & \-vma12\ & \-vma11\ & \-vma10\ & \-vma9\ & \-vma8\ & \-vma7\ & \-vma6\ & \-vma5\ & \-vma4\ & \-vma3\ & \-vma2\ & \-vma1\ & \-vma0\;
    \-md\ <= \-md31\ & \-md30\ & \-md29\ & \-md28\ & \-md27\ & \-md26\ & \-md25\ & \-md24\ & \-md23\ & \-md22\ & \-md21\ & \-md20\ & \-md19\ & \-md18\ & \-md17\ & \-md16\ & \-md15\ & \-md14\ & \-md13\ & \-md12\ & \-md11\ & \-md10\ & \-md9\ & \-md8\ & \-md7\ & \-md6\ & \-md5\ & \-md4\ & \-md3\ & \-md2\ & \-md1\ & \-md0\;
    alu <= alu32 & alu31 & alu30 & alu29 & alu28 & alu27 & alu26 & alu25 & alu24 & alu23 & alu22 & alu21 & alu20 & alu19 & alu18 & alu17 & alu16 & alu15 & alu14 & alu13 & alu12 & alu11 & alu10 & alu9 & alu8 & alu7 & alu6 & alu5 & alu4 & alu3 & alu2 & alu1 & alu0;
    q <= q31 & q30 & q29 & q28 & q27 & q26 & q25 & q24 & q23 & q22 & q21 & q20 & q19 & q18 & q17 & q16 & q15 & q14 & q13 & q12 & q11 & q10 & q9 & q8 & q7 & q6 & q5 & q4 & q3 & q2 & q1 & q0;
    r <= r31 & r30 & r29 & r28 & r27 & r26 & r25 & r24 & r23 & r22 & r21 & r20 & r19 & r18 & r17 & r16 & r15 & r14 & r13 & r12 & r11 & r10 & r9 & r8 & r7 & r6 & r5 & r4 & r3 & r2 & r1 & r0;
    aa <= aa17 & aa16 & aa15 & aa14 & aa13 & aa12 & aa11 & aa10 & aa9 & aa8 & aa7 & aa6 & aa5 & aa4 & aa3 & aa2 & aa1 & aa0;
    dc <= dc9 & dc8 & dc7 & dc6 & dc5 & dc4 & dc3 & dc2 & dc1 & dc0;
    dpc <= dpc13 & dpc12 & dpc11 & dpc10 & dpc9 & dpc8 & dpc7 & dpc6 & dpc5 & dpc4 & dpc3 & dpc2 & dpc1 & dpc0;
    iwr <= iwr48 & iwr47 & iwr46 & iwr45 & iwr44 & iwr43 & iwr42 & iwr41 & iwr40 & iwr39 & iwr38 & iwr37 & iwr36 & iwr35 & iwr34 & iwr33 & iwr32 & iwr31 & iwr30 & iwr29 & iwr28 & iwr27 & iwr26 & iwr25 & iwr24 & iwr23 & iwr22 & iwr21 & iwr20 & iwr19 & iwr18 & iwr17 & iwr16 & iwr15 & iwr14 & iwr13 & iwr12 & iwr11 & iwr10 & iwr9 & iwr8 & iwr7 & iwr6 & iwr5 & iwr4 & iwr3 & iwr2 & iwr1 & iwr0;
    lc <= lc25 & lc24 & lc23 & lc22 & lc21 & lc20 & lc19 & lc18 & lc17 & lc16 & lc15 & lc14 & lc13 & lc12 & lc11 & lc10 & lc9 & lc8 & lc7 & lc6 & lc5 & lc4 & lc3 & lc2 & lc1 & lc0;
    mapi <= mapi23 & mapi22 & mapi21 & mapi20 & mapi19 & mapi18 & mapi17 & mapi16 & mapi15 & mapi14 & mapi13 & mapi12 & mapi11 & mapi10 & mapi9 & mapi8;
    msk <= msk31 & msk30 & msk29 & msk28 & msk27 & msk26 & msk25 & msk24 & msk23 & msk22 & msk21 & msk20 & msk19 & msk18 & msk17 & msk16 & msk15 & msk14 & msk13 & msk12 & msk11 & msk10 & msk9 & msk8 & msk7 & msk6 & msk5 & msk4 & msk3 & msk2 & msk1 & msk0;
    opc <= opc13 & opc12 & opc11 & opc10 & opc9 & opc8 & opc7 & opc6 & opc5 & opc4 & opc3 & opc2 & opc1 & opc0;
    spc <= spc18 & spc17 & spc16 & spc15 & spc14 & spc13 & spc12 & spc11 & spc10 & spc9 & spc8 & spc7 & spc6 & spc5 & spc4 & spc3 & spc2 & spc1 & spc0;
    wadr <= wadr9 & wadr8 & wadr7 & wadr6 & wadr5 & wadr4 & wadr3 & wadr2 & wadr1 & wadr0;

    process (PC)
    begin
      if not is_x(PC) then
        if ((unsigned(PC) > 1) and (unsigned(PC) < 8#45#)) then
          report "PROM stucked at " & to_ostring(PC);
          std.env.stop;
        end if;
      end if;
    end process;

  end architecture;