library ieee;
use ieee.std_logic_1164.all;

package other is

end package other;

package body other is

end package body other;
