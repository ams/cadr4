library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity res20 is
  port (
    r2  : out std_logic; -- 2
    r3  : out std_logic; -- 3
    r4  : out std_logic; -- 4
    r5  : out std_logic; -- 5
    r6  : out std_logic; -- 6
    r7  : out std_logic; -- 7
    r8  : out std_logic; -- 8
    r9  : out std_logic; -- 9
    r10 : out std_logic; -- 10
    r11 : out std_logic; -- 11
    r12 : out std_logic; -- 12
    r13 : out std_logic; -- 13
    r14 : out std_logic; -- 14
    r15 : out std_logic; -- 15
    r16 : out std_logic; -- 16
    r17 : out std_logic; -- 17
    r18 : out std_logic; -- 18
    r19 : out std_logic -- 19
    );
end;

-- ChatGPT Codex implementation
architecture ttl of res20 is
begin
  r2  <= '1'; r3  <= '1'; r4  <= '1'; r5  <= '1';
  r6  <= '1'; r7  <= '1'; r8  <= '1'; r9  <= '1';
  r10 <= '1'; r11 <= '1'; r12 <= '1'; r13 <= '1';
  r14 <= '1'; r15 <= '1'; r16 <= '1'; r17 <= '1';
  r18 <= '1'; r19 <= '1';
end;
