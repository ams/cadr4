library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn7420_tb is
end sn7420_tb;

architecture testbench of sn7420_tb is

begin

--  uut : sn7420 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
