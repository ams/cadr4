library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_vmemdr is
  port (
    \-mapdrive\ : out std_logic;
    \-pfw\      : in  std_logic;
    mf24        : out std_logic;
    \-pfr\      : in  std_logic;
    mf25        : out std_logic;
    hi12        : in  std_logic;
    mf26        : out std_logic;
    \-vmap4\    : in  std_logic;
    mf27        : out std_logic;
    \-vmap3\    : in  std_logic;
    mf28        : out std_logic;
    \-vmap2\    : in  std_logic;
    mf29        : out std_logic;
    \-vmap1\    : in  std_logic;
    mf30        : out std_logic;
    \-vmap0\    : in  std_logic;
    mf31        : out std_logic;
    \-vmo15\    : in  std_logic;
    mf8         : out std_logic;
    \-vmo14\    : in  std_logic;
    mf9         : out std_logic;
    \-vmo13\    : in  std_logic;
    mf10        : out std_logic;
    \-vmo12\    : in  std_logic;
    mf11        : out std_logic;
    \-vmo11\    : in  std_logic;
    mf12        : out std_logic;
    \-vmo10\    : in  std_logic;
    mf13        : out std_logic;
    \-vmo9\     : in  std_logic;
    mf14        : out std_logic;
    \-vmo8\     : in  std_logic;
    mf15        : out std_logic;
    \-vmo23\    : in  std_logic;
    mf16        : out std_logic;
    \-vmo22\    : in  std_logic;
    mf17        : out std_logic;
    \-vmo21\    : in  std_logic;
    mf18        : out std_logic;
    \-vmo20\    : in  std_logic;
    mf19        : out std_logic;
    \-vmo19\    : in  std_logic;
    mf20        : out std_logic;
    \-vmo18\    : in  std_logic;
    mf21        : out std_logic;
    \-vmo17\    : in  std_logic;
    mf22        : out std_logic;
    \-vmo16\    : in  std_logic;
    mf23        : out std_logic;
    tse1a       : in  std_logic;
    srcmap      : out std_logic;
    \-vmo7\     : in  std_logic;
    mf0         : out std_logic;
    \-vmo6\     : in  std_logic;
    mf1         : out std_logic;
    \-vmo5\     : in  std_logic;
    mf2         : out std_logic;
    \-vmo4\     : in  std_logic;
    mf3         : out std_logic;
    \-vmo3\     : in  std_logic;
    mf4         : out std_logic;
    \-vmo2\     : in  std_logic;
    mf5         : out std_logic;
    \-vmo1\     : in  std_logic;
    mf6         : out std_logic;
    \-vmo0\     : in  std_logic;
    mf7         : out std_logic;
    gnd         : in  std_logic;
    \-lvmo23\   : out std_logic;
    \-lvmo22\   : out std_logic;
    \-pma21\    : out std_logic;
    \-pma20\    : out std_logic;
    memstart    : in  std_logic;
    \-pma19\    : out std_logic;
    \-pma18\    : out std_logic;
    \-pma17\    : out std_logic;
    \-pma16\    : out std_logic;
    \-pma15\    : out std_logic;
    \-pma14\    : out std_logic;
    \-pma13\    : out std_logic;
    \-pma12\    : out std_logic;
    \-pma11\    : out std_logic;
    \-pma10\    : out std_logic;
    \-pma9\     : out std_logic;
    \-pma8\     : out std_logic;
    \-vma6\     : in  std_logic;
    \-vma5\     : in  std_logic;
    \-vma4\     : in  std_logic;
    \-vma3\     : in  std_logic;
    \-vma2\     : in  std_logic;
    \-vma1\     : in  std_logic;
    \-vma0\     : in  std_logic;
    \-vma7\     : in  std_logic;
    \-adrpar\   : out std_logic;
    \-srcmap\   : in  std_logic);
end;

architecture ttl of cadr4_vmemdr is
  signal internal13 : std_logic;
  signal nc100      : std_logic;
  signal nc99       : std_logic;
begin
  vmemdr_1a01 : sn74s240 port map(aenb_n => \-mapdrive\, ain0 => \-pfw\, bout3 => mf24, ain1 => \-pfr\, bout2 => mf25, ain2 => hi12, bout1 => mf26, ain3 => \-vmap4\, bout0 => mf27, bin0 => \-vmap3\, aout3 => mf28, bin1 => \-vmap2\, aout2 => mf29, bin2 => \-vmap1\, aout1 => mf30, bin3 => \-vmap0\, aout0 => mf31, benb_n => \-mapdrive\);
  vmemdr_1a03 : sn74s240 port map(aenb_n => \-mapdrive\, ain0 => \-vmo15\, bout3 => mf8, ain1 => \-vmo14\, bout2 => mf9, ain2 => \-vmo13\, bout1 => mf10, ain3 => \-vmo12\, bout0 => mf11, bin0 => \-vmo11\, aout3 => mf12, bin1 => \-vmo10\, aout2 => mf13, bin2 => \-vmo9\, aout1 => mf14, bin3 => \-vmo8\, aout0 => mf15, benb_n => \-mapdrive\);
  vmemdr_1a07 : sn74s240 port map(aenb_n => \-mapdrive\, ain0 => \-vmo23\, bout3 => mf16, ain1 => \-vmo22\, bout2 => mf17, ain2 => \-vmo21\, bout1 => mf18, ain3 => \-vmo20\, bout0 => mf19, bin0 => \-vmo19\, aout3 => mf20, bin1 => \-vmo18\, aout2 => mf21, bin2 => \-vmo17\, aout1 => mf22, bin3 => \-vmo16\, aout0 => mf23, benb_n => \-mapdrive\);
  vmemdr_1a08 : sn74s00 port map(g1b     => tse1a, g1a => srcmap, g1q_n => \-mapdrive\, g2b => '0', g2a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  vmemdr_1a13 : sn74s240 port map(aenb_n => \-mapdrive\, ain0 => \-vmo7\, bout3 => mf0, ain1 => \-vmo6\, bout2 => mf1, ain2 => \-vmo5\, bout1 => mf2, ain3 => \-vmo4\, bout0 => mf3, bin0 => \-vmo3\, aout3 => mf4, bin1 => \-vmo2\, aout2 => mf5, bin2 => \-vmo1\, aout1 => mf6, bin3 => \-vmo0\, aout0 => mf7, benb_n => \-mapdrive\);
  vmemdr_1d14 : sn74s373 port map(oenb_n => gnd, o0 => \-lvmo23\, i0 => \-vmo23\, i1 => \-vmo22\, o1 => \-lvmo22\, o2 => \-pma21\, i2 => \-vmo13\, i3 => \-vmo12\, o3 => \-pma20\, hold_n => memstart, o4 => \-pma19\, i4 => \-vmo11\, i5 => \-vmo10\, o5 => \-pma18\, o6 => \-pma17\, i6 => \-vmo9\, i7 => \-vmo8\, o7 => \-pma16\);
  vmemdr_1d15 : sn74s373 port map(oenb_n => gnd, o0 => \-pma15\, i0 => \-vmo7\, i1 => \-vmo6\, o1 => \-pma14\, o2 => \-pma13\, i2 => \-vmo5\, i3 => \-vmo4\, o3 => \-pma12\, hold_n => memstart, o4 => \-pma11\, i4 => \-vmo3\, i5 => \-vmo2\, o5 => \-pma10\, o6 => \-pma9\, i6 => \-vmo1\, i7 => \-vmo0\, o7 => \-pma8\);
  vmemdr_1e17 : am93s48 port map(i6      => \-vma6\, i5 => \-vma5\, i4 => \-vma4\, i3 => \-vma3\, i2 => \-vma2\, i1 => \-vma1\, i0 => \-vma0\, po => internal13, pe => nc100, i11 => \-pma11\, i10 => \-pma10\, i9 => \-pma9\, i8 => \-pma8\, i7 => \-vma7\);
  vmemdr_1e18 : am93s48 port map(i6      => \-pma18\, i5 => \-pma17\, i4 => \-pma16\, i3 => \-pma15\, i2 => \-pma14\, i1 => \-pma13\, i0 => \-pma12\, po => \-adrpar\, pe => nc99, i11 => internal13, i10 => gnd, i9 => \-pma21\, i8 => \-pma20\, i7 => \-pma19\);
  vmemdr_2a05 : sn74s04 port map(g4q_n   => srcmap, g4a => \-srcmap\, g1a => '0', g2a => '0', g3a => '0', g5a => '0', g6a => '0');
end architecture;
