library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_spy1 is
  port (
    \-spy.obl\ : out std_logic;
    ob7        : in  std_logic;
    spy0       : out std_logic;
    ob6        : in  std_logic;
    spy1       : out std_logic;
    ob5        : in  std_logic;
    spy2       : out std_logic;
    ob4        : in  std_logic;
    spy3       : out std_logic;
    ob3        : in  std_logic;
    spy4       : out std_logic;
    ob2        : in  std_logic;
    spy5       : out std_logic;
    ob1        : in  std_logic;
    spy6       : out std_logic;
    ob0        : in  std_logic;
    spy7       : out std_logic;
    ob15       : in  std_logic;
    spy8       : out std_logic;
    ob14       : in  std_logic;
    spy9       : out std_logic;
    ob13       : in  std_logic;
    spy10      : out std_logic;
    ob12       : in  std_logic;
    spy11      : out std_logic;
    ob11       : in  std_logic;
    spy12      : out std_logic;
    ob10       : in  std_logic;
    spy13      : out std_logic;
    ob9        : in  std_logic;
    spy14      : out std_logic;
    ob8        : in  std_logic;
    spy15      : out std_logic;
    \-spy.obh\ : in  std_logic;
    ob23       : in  std_logic;
    ob22       : in  std_logic;
    ob21       : in  std_logic;
    ob20       : in  std_logic;
    ob19       : in  std_logic;
    ob18       : in  std_logic;
    ob17       : in  std_logic;
    ob16       : in  std_logic;
    ob31       : in  std_logic;
    ob30       : in  std_logic;
    ob29       : in  std_logic;
    ob28       : in  std_logic;
    ob27       : in  std_logic;
    ob26       : in  std_logic;
    ob25       : in  std_logic;
    ob24       : in  std_logic;
    \-spy.irl\ : in  std_logic;
    ir7        : in  std_logic;
    ir6        : in  std_logic;
    ir5        : in  std_logic;
    ir4        : in  std_logic;
    ir3        : in  std_logic;
    ir2        : in  std_logic;
    ir1        : in  std_logic;
    ir0        : in  std_logic;
    ir15       : in  std_logic;
    ir14       : in  std_logic;
    ir13       : in  std_logic;
    ir12       : in  std_logic;
    ir11       : in  std_logic;
    ir10       : in  std_logic;
    ir9        : in  std_logic;
    ir8        : in  std_logic;
    \-spy.irh\ : in  std_logic;
    ir47       : in  std_logic;
    ir46       : in  std_logic;
    ir45       : in  std_logic;
    ir44       : in  std_logic;
    ir43       : in  std_logic;
    ir42       : in  std_logic;
    ir41       : in  std_logic;
    ir40       : in  std_logic;
    ir39       : in  std_logic;
    ir38       : in  std_logic;
    ir37       : in  std_logic;
    ir36       : in  std_logic;
    ir35       : in  std_logic;
    ir34       : in  std_logic;
    ir33       : in  std_logic;
    ir32       : in  std_logic;
    \-spy.irm\ : in  std_logic;
    ir31       : in  std_logic;
    ir30       : in  std_logic;
    ir29       : in  std_logic;
    ir28       : in  std_logic;
    ir27       : in  std_logic;
    ir26       : in  std_logic;
    ir25       : in  std_logic;
    ir24       : in  std_logic;
    ir23       : in  std_logic;
    ir22       : in  std_logic;
    ir21       : in  std_logic;
    ir20       : in  std_logic;
    ir19       : in  std_logic;
    ir18       : in  std_logic;
    ir17       : in  std_logic;
    ir16       : in  std_logic);
end;

architecture ttl of cadr4_spy1 is
begin
  spy1_2c17 : sn74ls244 port map(aenb_n => \-spy.obl\, ain0 => ob7, bout3 => spy0, ain1 => ob6, bout2 => spy1, ain2 => ob5, bout1 => spy2, ain3 => ob4, bout0 => spy3, bin0 => ob3, aout3 => spy4, bin1 => ob2, aout2 => spy5, bin2 => ob1, aout1 => spy6, bin3 => ob0, aout0 => spy7, benb_n => \-spy.obl\);
  spy1_2c18 : sn74ls244 port map(aenb_n => \-spy.obl\, ain0 => ob15, bout3 => spy8, ain1 => ob14, bout2 => spy9, ain2 => ob13, bout1 => spy10, ain3 => ob12, bout0 => spy11, bin0 => ob11, aout3 => spy12, bin1 => ob10, aout2 => spy13, bin2 => ob9, aout1 => spy14, bin3 => ob8, aout0 => spy15, benb_n => \-spy.obl\);
  spy1_3c23 : sn74ls244 port map(aenb_n => \-spy.obh\, ain0 => ob23, bout3 => spy0, ain1 => ob22, bout2 => spy1, ain2 => ob21, bout1 => spy2, ain3 => ob20, bout0 => spy3, bin0 => ob19, aout3 => spy4, bin1 => ob18, aout2 => spy5, bin2 => ob17, aout1 => spy6, bin3 => ob16, aout0 => spy7, benb_n => \-spy.obh\);
  spy1_3c24 : sn74ls244 port map(aenb_n => \-spy.obh\, ain0 => ob31, bout3 => spy8, ain1 => ob30, bout2 => spy9, ain2 => ob29, bout1 => spy10, ain3 => ob28, bout0 => spy11, bin0 => ob27, aout3 => spy12, bin1 => ob26, aout2 => spy13, bin2 => ob25, aout1 => spy14, bin3 => ob24, aout0 => spy15, benb_n => \-spy.obh\);
  spy1_3e01 : sn74ls244 port map(aenb_n => \-spy.irl\, ain0 => ir7, bout3 => spy0, ain1 => ir6, bout2 => spy1, ain2 => ir5, bout1 => spy2, ain3 => ir4, bout0 => spy3, bin0 => ir3, aout3 => spy4, bin1 => ir2, aout2 => spy5, bin2 => ir1, aout1 => spy6, bin3 => ir0, aout0 => spy7, benb_n => \-spy.irl\);
  spy1_3e03 : sn74ls244 port map(aenb_n => \-spy.irl\, ain0 => ir15, bout3 => spy8, ain1 => ir14, bout2 => spy9, ain2 => ir13, bout1 => spy10, ain3 => ir12, bout0 => spy11, bin0 => ir11, aout3 => spy12, bin1 => ir10, aout2 => spy13, bin2 => ir9, aout1 => spy14, bin3 => ir8, aout0 => spy15, benb_n => \-spy.irl\);
  spy1_3e06 : sn74ls244 port map(aenb_n => \-spy.irh\, ain0 => ir47, bout3 => spy8, ain1 => ir46, bout2 => spy9, ain2 => ir45, bout1 => spy10, ain3 => ir44, bout0 => spy11, bin0 => ir43, aout3 => spy12, bin1 => ir42, aout2 => spy13, bin2 => ir41, aout1 => spy14, bin3 => ir40, aout0 => spy15, benb_n => \-spy.irh\);
  spy1_3f21 : sn74ls244 port map(aenb_n => \-spy.irh\, ain0 => ir39, bout3 => spy0, ain1 => ir38, bout2 => spy1, ain2 => ir37, bout1 => spy2, ain3 => ir36, bout0 => spy3, bin0 => ir35, aout3 => spy4, bin1 => ir34, aout2 => spy5, bin2 => ir33, aout1 => spy6, bin3 => ir32, aout0 => spy7, benb_n => \-spy.irh\);
  spy1_3f23 : sn74ls244 port map(aenb_n => \-spy.irm\, ain0 => ir31, bout3 => spy8, ain1 => ir30, bout2 => spy9, ain2 => ir29, bout1 => spy10, ain3 => ir28, bout0 => spy11, bin0 => ir27, aout3 => spy12, bin1 => ir26, aout2 => spy13, bin2 => ir25, aout1 => spy14, bin3 => ir24, aout0 => spy15, benb_n => \-spy.irm\);
  spy1_3f25 : sn74ls244 port map(aenb_n => \-spy.irm\, ain0 => ir23, bout3 => spy0, ain1 => ir22, bout2 => spy1, ain2 => ir21, bout1 => spy2, ain3 => ir20, bout0 => spy3, bin0 => ir19, aout3 => spy4, bin1 => ir18, aout2 => spy5, bin2 => ir17, aout1 => spy6, bin3 => ir16, aout0 => spy7, benb_n => \-spy.irm\);
end architecture;
