library ieee;
use ieee.std_logic_1164.all;

entity ic_16dummy_tb is
end;

architecture testbench of ic_16dummy_tb is

  signal \-boot2\       : std_logic;
  signal \-power reset\ : std_logic;

begin

  uut : entity work.ic_16dummy port map(
    \-boot2\ => \-boot2\,
    \-power reset\ => \-power reset\
    );

  process
  begin
    -- Test static outputs
    assert \-boot2\ = 'H' report "-boot2 should be 'H'";
    assert \-power reset\ = '0' report "-power reset should be '0' initially";
    wait for 20 ns;
    assert \-power reset\ = '1' report "-power reset should be '1' after delay";
    wait;
  end process;

end;
