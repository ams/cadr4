library ieee;
use ieee.std_logic_1164.all;

entity busint_uprior is
  port (
    \-clk\          : in     std_logic;
    \-disable int grant\ : in     std_logic;
    \-local enable\ : in     std_logic;
    \-npg out\      : in     std_logic;
    \bus req\       : in     std_logic;
    \local enable\  : in     std_logic;
    \sack in\       : in     std_logic;
    level0          : in     std_logic;
    level1          : in     std_logic;
    reset           : in     std_logic;
    \-ub br4\       : inout  std_logic;
    \-ub br5\       : inout  std_logic;
    \-ub br6\       : inout  std_logic;
    \-ub br7\       : inout  std_logic;
    \-ub init\      : inout  std_logic;
    \-ub intr\      : inout  std_logic;
    \-ub npr\       : inout  std_logic;
    \hi 1-14\       : inout  std_logic;
    \ub npg in\     : inout  std_logic;
    \ub npg out\    : inout  std_logic;
    \-any grant dlyd\ : out    std_logic;
    \-bg4o\         : out    std_logic;
    \-bg5o\         : out    std_logic;
    \-bg6o\         : out    std_logic;
    \-bg7o\         : out    std_logic;
    \-clear grant\  : out    std_logic;
    \-npg in\       : out    std_logic;
    \-npgo\         : out    std_logic;
    \any grant dlyd\ : out    std_logic;
    \any grant\     : out    std_logic;
    \any int grant\ : out    std_logic;
    \grant timeout\ : out    std_logic;
    \ub bg4 in\     : out    std_logic;
    \ub bg5 in\     : out    std_logic;
    \ub bg6 in\     : out    std_logic;
    \ub bg7 in\     : out    std_logic;
    \unibus init in\ : out    std_logic;
    \unibus intr in\ : out    std_logic;
    bg4o            : out    std_logic;
    bg4p            : out    std_logic;
    bg5o            : out    std_logic;
    bg5p            : out    std_logic;
    bg6o            : out    std_logic;
    bg6p            : out    std_logic;
    bg7o            : out    std_logic;
    bg7p            : out    std_logic;
    br4             : out    std_logic;
    br4d            : out    std_logic;
    br5             : out    std_logic;
    br5d            : out    std_logic;
    br6             : out    std_logic;
    br6d            : out    std_logic;
    br7             : out    std_logic;
    br7d            : out    std_logic;
    npgo            : out    std_logic;
    npgp            : out    std_logic;
    npr             : out    std_logic;
    nprd            : out    std_logic;
    sackd           : out    std_logic
  );
end entity;
