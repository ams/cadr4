library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_mmem is
  port (
    \-mwpa\    : in  std_logic;
    gnd        : in  std_logic;
    l16        : in  std_logic;
    \-madr4a\  : in  std_logic;
    hi3        : in  std_logic;
    mmem16     : out std_logic;
    mmem17     : out std_logic;
    \-madr3a\  : in  std_logic;
    \-madr2a\  : in  std_logic;
    \-madr1a\  : in  std_logic;
    \-madr0a\  : in  std_logic;
    l17        : in  std_logic;
    \-mwpb\    : in  std_logic;
    l12        : in  std_logic;
    \-madr4b\  : in  std_logic;
    hi2        : in  std_logic;
    mmem12     : out std_logic;
    mmem13     : out std_logic;
    \-madr3b\  : in  std_logic;
    \-madr2b\  : in  std_logic;
    \-madr1b\  : in  std_logic;
    \-madr0b\  : in  std_logic;
    l13        : in  std_logic;
    l8         : in  std_logic;
    mmem8      : out std_logic;
    mmem9      : out std_logic;
    l9         : in  std_logic;
    l4         : in  std_logic;
    mmem4      : out std_logic;
    mmem5      : out std_logic;
    l5         : in  std_logic;
    l0         : in  std_logic;
    mmem0      : out std_logic;
    mmem1      : out std_logic;
    l1         : in  std_logic;
    l18        : in  std_logic;
    mmem18     : out std_logic;
    mmem19     : out std_logic;
    l19        : in  std_logic;
    l14        : in  std_logic;
    mmem14     : out std_logic;
    mmem15     : out std_logic;
    l15        : in  std_logic;
    l10        : in  std_logic;
    mmem10     : out std_logic;
    mmem11     : out std_logic;
    l11        : in  std_logic;
    l6         : in  std_logic;
    mmem6      : out std_logic;
    mmem7      : out std_logic;
    l7         : in  std_logic;
    l2         : in  std_logic;
    mmem2      : out std_logic;
    mmem3      : out std_logic;
    l3         : in  std_logic;
    l28        : in  std_logic;
    mmem28     : out std_logic;
    mmem29     : out std_logic;
    l29        : in  std_logic;
    l24        : in  std_logic;
    mmem24     : out std_logic;
    mmem25     : out std_logic;
    l25        : in  std_logic;
    l20        : in  std_logic;
    mmem20     : out std_logic;
    mmem21     : out std_logic;
    l21        : in  std_logic;
    lparity    : in  std_logic;
    mmemparity : out std_logic;
    l30        : in  std_logic;
    mmem30     : out std_logic;
    mmem31     : out std_logic;
    l31        : in  std_logic;
    l26        : in  std_logic;
    mmem26     : out std_logic;
    mmem27     : out std_logic;
    l27        : in  std_logic;
    l22        : in  std_logic;
    mmem22     : out std_logic;
    mmem23     : out std_logic;
    l23        : in  std_logic);
end;

architecture ttl of cadr_mmem is
  signal nc291 : std_logic;
  signal nc292 : std_logic;
  signal nc293 : std_logic;
begin
  mmem_4a21 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l16, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem16, d1 => mmem17, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l17, we1_n => gnd);
  mmem_4a22 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l12, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem12, d1 => mmem13, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l13, we1_n => gnd);
  mmem_4a23 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l8, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem8, d1 => mmem9, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l9, we1_n => gnd);
  mmem_4a24 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l4, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem4, d1 => mmem5, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l5, we1_n => gnd);
  mmem_4a25 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l0, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem0, d1 => mmem1, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l1, we1_n => gnd);
  mmem_4a26 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l18, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem18, d1 => mmem19, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l19, we1_n => gnd);
  mmem_4a27 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l14, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem14, d1 => mmem15, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l15, we1_n => gnd);
  mmem_4a28 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l10, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem10, d1 => mmem11, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l11, we1_n => gnd);
  mmem_4a29 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l6, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem6, d1 => mmem7, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l7, we1_n => gnd);
  mmem_4a30 : dm82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l2, a4 => \-madr4b\, ce => hi2, strobe => hi2, d0 => mmem2, d1 => mmem3, a3 => \-madr3b\, a2 => \-madr2b\, a1 => \-madr1b\, a0 => \-madr0b\, i1 => l3, we1_n => gnd);
  mmem_4b23 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l28, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem28, d1 => mmem29, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l29, we1_n => gnd);
  mmem_4b24 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l24, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem24, d1 => mmem25, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l25, we1_n => gnd);
  mmem_4b25 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l20, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem20, d1 => mmem21, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l21, we1_n => gnd);
  mmem_4b27 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => lparity, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmemparity, d1 => nc291, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => nc292, we1_n => nc293);
  mmem_4b28 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l30, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem30, d1 => mmem31, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l31, we1_n => gnd);
  mmem_4b29 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l26, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem26, d1 => mmem27, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l27, we1_n => gnd);
  mmem_4b30 : dm82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l22, a4 => \-madr4a\, ce => hi3, strobe => hi3, d0 => mmem22, d1 => mmem23, a3 => \-madr3a\, a2 => \-madr2a\, a1 => \-madr1a\, a0 => \-madr0a\, i1 => l23, we1_n => gnd);
end architecture;
