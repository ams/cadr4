library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_mo0 is
  port (
    alu15  : in  std_logic;
    r15    : in  std_logic;
    a15    : in  std_logic;
    ob15   : out std_logic;
    gnd    : in  std_logic;
    osel1b : in  std_logic;
    osel0b : in  std_logic;
    msk15  : in  std_logic;
    alu14  : in  std_logic;
    alu16  : in  std_logic;
    r14    : in  std_logic;
    a14    : in  std_logic;
    ob14   : out std_logic;
    msk14  : in  std_logic;
    alu13  : in  std_logic;
    r13    : in  std_logic;
    a13    : in  std_logic;
    ob13   : out std_logic;
    msk13  : in  std_logic;
    alu12  : in  std_logic;
    r12    : in  std_logic;
    a12    : in  std_logic;
    ob12   : out std_logic;
    msk12  : in  std_logic;
    alu11  : in  std_logic;
    alu7   : in  std_logic;
    r7     : in  std_logic;
    a7     : in  std_logic;
    ob7    : out std_logic;
    msk7   : in  std_logic;
    alu6   : in  std_logic;
    alu8   : in  std_logic;
    r6     : in  std_logic;
    a6     : in  std_logic;
    ob6    : out std_logic;
    msk6   : in  std_logic;
    alu5   : in  std_logic;
    r5     : in  std_logic;
    a5     : in  std_logic;
    ob5    : out std_logic;
    msk5   : in  std_logic;
    alu4   : in  std_logic;
    r4     : in  std_logic;
    a4     : in  std_logic;
    ob4    : out std_logic;
    msk4   : in  std_logic;
    alu3   : in  std_logic;
    r11    : in  std_logic;
    a11    : in  std_logic;
    ob11   : out std_logic;
    msk11  : in  std_logic;
    alu10  : in  std_logic;
    r10    : in  std_logic;
    a10    : in  std_logic;
    ob10   : out std_logic;
    msk10  : in  std_logic;
    alu9   : in  std_logic;
    r3     : in  std_logic;
    a3     : in  std_logic;
    ob3    : out std_logic;
    msk3   : in  std_logic;
    alu2   : in  std_logic;
    r2     : in  std_logic;
    a2     : in  std_logic;
    ob2    : out std_logic;
    msk2   : in  std_logic;
    alu1   : in  std_logic;
    r9     : in  std_logic;
    a9     : in  std_logic;
    ob9    : out std_logic;
    msk9   : in  std_logic;
    r8     : in  std_logic;
    a8     : in  std_logic;
    ob8    : out std_logic;
    msk8   : in  std_logic;
    r1     : in  std_logic;
    a1     : in  std_logic;
    ob1    : out std_logic;
    msk1   : in  std_logic;
    alu0   : in  std_logic;
    r0     : in  std_logic;
    a0     : in  std_logic;
    ob0    : out std_logic;
    msk0   : in  std_logic;
    q31    : in  std_logic);
end;

architecture ttl of cadr4_mo0 is
  signal nc275 : std_logic;
  signal nc276 : std_logic;
  signal nc277 : std_logic;
  signal nc278 : std_logic;
  signal nc279 : std_logic;
  signal nc280 : std_logic;
  signal nc281 : std_logic;
  signal nc282 : std_logic;
  signal nc283 : std_logic;
  signal nc284 : std_logic;
  signal nc285 : std_logic;
  signal nc286 : std_logic;
  signal nc287 : std_logic;
  signal nc288 : std_logic;
  signal nc289 : std_logic;
  signal nc290 : std_logic;
begin
  mo0_2a24 : sn74s151 port map(i3 => alu15, i2 => alu15, i1 => r15, i0 => a15, q => ob15, q_n => nc290, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk15, i7 => alu14, i6 => alu14, i5 => alu16, i4 => alu16);
  mo0_2a25 : sn74s151 port map(i3 => alu14, i2 => alu14, i1 => r14, i0 => a14, q => ob14, q_n => nc289, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk14, i7 => alu13, i6 => alu13, i5 => alu15, i4 => alu15);
  mo0_2a29 : sn74s151 port map(i3 => alu13, i2 => alu13, i1 => r13, i0 => a13, q => ob13, q_n => nc288, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk13, i7 => alu12, i6 => alu12, i5 => alu14, i4 => alu14);
  mo0_2a30 : sn74s151 port map(i3 => alu12, i2 => alu12, i1 => r12, i0 => a12, q => ob12, q_n => nc287, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk12, i7 => alu11, i6 => alu11, i5 => alu13, i4 => alu13);
  mo0_2b24 : sn74s151 port map(i3 => alu7, i2 => alu7, i1 => r7, i0 => a7, q => ob7, q_n => nc282, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk7, i7 => alu6, i6 => alu6, i5 => alu8, i4 => alu8);
  mo0_2b25 : sn74s151 port map(i3 => alu6, i2 => alu6, i1 => r6, i0 => a6, q => ob6, q_n => nc281, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk6, i7 => alu5, i6 => alu5, i5 => alu7, i4 => alu7);
  mo0_2b29 : sn74s151 port map(i3 => alu5, i2 => alu5, i1 => r5, i0 => a5, q => ob5, q_n => nc280, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk5, i7 => alu4, i6 => alu4, i5 => alu6, i4 => alu6);
  mo0_2b30 : sn74s151 port map(i3 => alu4, i2 => alu4, i1 => r4, i0 => a4, q => ob4, q_n => nc279, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk4, i7 => alu3, i6 => alu3, i5 => alu5, i4 => alu5);
  mo0_2c19 : sn74s151 port map(i3 => alu11, i2 => alu11, i1 => r11, i0 => a11, q => ob11, q_n => nc286, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk11, i7 => alu10, i6 => alu10, i5 => alu12, i4 => alu12);
  mo0_2c24 : sn74s151 port map(i3 => alu10, i2 => alu10, i1 => r10, i0 => a10, q => ob10, q_n => nc285, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk10, i7 => alu9, i6 => alu9, i5 => alu11, i4 => alu11);
  mo0_2c29 : sn74s151 port map(i3 => alu3, i2 => alu3, i1 => r3, i0 => a3, q => ob3, q_n => nc278, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk3, i7 => alu2, i6 => alu2, i5 => alu4, i4 => alu4);
  mo0_2c30 : sn74s151 port map(i3 => alu2, i2 => alu2, i1 => r2, i0 => a2, q => ob2, q_n => nc277, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk2, i7 => alu1, i6 => alu1, i5 => alu3, i4 => alu3);
  mo0_2d23 : sn74s151 port map(i3 => alu9, i2 => alu9, i1 => r9, i0 => a9, q => ob9, q_n => nc284, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk9, i7 => alu8, i6 => alu8, i5 => alu10, i4 => alu10);
  mo0_2d24 : sn74s151 port map(i3 => alu8, i2 => alu8, i1 => r8, i0 => a8, q => ob8, q_n => nc283, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk8, i7 => alu7, i6 => alu7, i5 => alu9, i4 => alu9);
  mo0_2d28 : sn74s151 port map(i3 => alu1, i2 => alu1, i1 => r1, i0 => a1, q => ob1, q_n => nc276, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk1, i7 => alu0, i6 => alu0, i5 => alu2, i4 => alu2);
  mo0_2d29 : sn74s151 port map(i3 => alu0, i2 => alu0, i1 => r0, i0 => a0, q => ob0, q_n => nc275, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk0, i7 => q31, i6 => q31, i5 => alu1, i4 => alu1);
end architecture;
