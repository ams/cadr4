library ieee;
use ieee.std_logic_1164.all;

entity icmem_iram31 is
  port (
    \-ice1d\        : in     std_logic;
    \-iwen\         : in     std_logic;
    \-pcc0\         : in     std_logic;
    \-pcc10\        : in     std_logic;
    \-pcc11\        : in     std_logic;
    \-pcc1\         : in     std_logic;
    \-pcc2\         : in     std_logic;
    \-pcc3\         : in     std_logic;
    \-pcc4\         : in     std_logic;
    \-pcc5\         : in     std_logic;
    \-pcc6\         : in     std_logic;
    \-pcc7\         : in     std_logic;
    \-pcc8\         : in     std_logic;
    \-pcc9\         : in     std_logic;
    iwr36           : in     std_logic;
    iwr37           : in     std_logic;
    iwr38           : in     std_logic;
    iwr39           : in     std_logic;
    iwr40           : in     std_logic;
    iwr41           : in     std_logic;
    iwr42           : in     std_logic;
    iwr43           : in     std_logic;
    iwr44           : in     std_logic;
    iwr45           : in     std_logic;
    iwr46           : in     std_logic;
    iwr47           : in     std_logic;
    iwr48           : in     std_logic;
    i36             : out    std_logic;
    i37             : out    std_logic;
    i38             : out    std_logic;
    i39             : out    std_logic;
    i40             : out    std_logic;
    i41             : out    std_logic;
    i42             : out    std_logic;
    i43             : out    std_logic;
    i44             : out    std_logic;
    i45             : out    std_logic;
    i46             : out    std_logic;
    i47             : out    std_logic;
    i48             : out    std_logic;
    pc0n            : out    std_logic;
    pc10n           : out    std_logic;
    pc11n           : out    std_logic;
    pc1n            : out    std_logic;
    pc2n            : out    std_logic;
    pc3n            : out    std_logic;
    pc4n            : out    std_logic;
    pc5n            : out    std_logic;
    pc6n            : out    std_logic;
    pc7n            : out    std_logic;
    pc8n            : out    std_logic;
    pc9n            : out    std_logic
  );
end entity;
