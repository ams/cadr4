library ieee;
use ieee.std_logic_1164.all;

entity cadr_dspctl is
  port (
    \-funct2\       : in     std_logic;
    \-irdisp\       : in     std_logic;
    a0              : in     std_logic;
    a1              : in     std_logic;
    a10             : in     std_logic;
    a11             : in     std_logic;
    a12             : in     std_logic;
    a13             : in     std_logic;
    a14             : in     std_logic;
    a15             : in     std_logic;
    a16             : in     std_logic;
    a17             : in     std_logic;
    a2              : in     std_logic;
    a3              : in     std_logic;
    a4              : in     std_logic;
    a5              : in     std_logic;
    a6              : in     std_logic;
    a7              : in     std_logic;
    a8              : in     std_logic;
    a9              : in     std_logic;
    clk3e           : in     std_logic;
    dispenb         : in     std_logic;
    dn              : in     std_logic;
    dp              : in     std_logic;
    dpar            : in     std_logic;
    dpc0            : in     std_logic;
    dpc1            : in     std_logic;
    dpc10           : in     std_logic;
    dpc11           : in     std_logic;
    dpc12           : in     std_logic;
    dpc13           : in     std_logic;
    dpc2            : in     std_logic;
    dpc3            : in     std_logic;
    dpc4            : in     std_logic;
    dpc5            : in     std_logic;
    dpc6            : in     std_logic;
    dpc7            : in     std_logic;
    dpc8            : in     std_logic;
    dpc9            : in     std_logic;
    dr              : in     std_logic;
    hi4             : in     std_logic;
    ir32            : in     std_logic;
    ir33            : in     std_logic;
    ir34            : in     std_logic;
    ir35            : in     std_logic;
    ir36            : in     std_logic;
    ir37            : in     std_logic;
    ir38            : in     std_logic;
    ir39            : in     std_logic;
    ir40            : in     std_logic;
    ir41            : in     std_logic;
    ir5             : in     std_logic;
    ir6             : in     std_logic;
    ir7             : in     std_logic;
    ir8             : in     std_logic;
    ir9             : in     std_logic;
    \-dmapbenb\     : out    std_logic;
    \-dparh\        : out    std_logic;
    aa0             : out    std_logic;
    aa1             : out    std_logic;
    aa10            : out    std_logic;
    aa11            : out    std_logic;
    aa12            : out    std_logic;
    aa13            : out    std_logic;
    aa14            : out    std_logic;
    aa15            : out    std_logic;
    aa16            : out    std_logic;
    aa17            : out    std_logic;
    aa2             : out    std_logic;
    aa3             : out    std_logic;
    aa4             : out    std_logic;
    aa5             : out    std_logic;
    aa6             : out    std_logic;
    aa7             : out    std_logic;
    aa8             : out    std_logic;
    aa9             : out    std_logic;
    dc0             : out    std_logic;
    dc1             : out    std_logic;
    dc2             : out    std_logic;
    dc3             : out    std_logic;
    dc4             : out    std_logic;
    dc5             : out    std_logic;
    dc6             : out    std_logic;
    dc7             : out    std_logic;
    dc8             : out    std_logic;
    dc9             : out    std_logic;
    dispwr          : out    std_logic;
    dmask0          : out    std_logic;
    dmask1          : out    std_logic;
    dmask2          : out    std_logic;
    dmask3          : out    std_logic;
    dmask4          : out    std_logic;
    dmask5          : out    std_logic;
    dmask6          : out    std_logic;
    dpareven        : out    std_logic;
    dparl           : out    std_logic;
    dparok          : out    std_logic
  );
end entity cadr_dspctl;
