library ieee;
use ieee.std_logic_1164.all;

entity cadr_pdl1 is
  port (
    \-pdla0a\ : in  std_logic;
    \-pdla1a\ : in  std_logic;
    \-pdla2a\ : in  std_logic;
    \-pdla3a\ : in  std_logic;
    \-pdla4a\ : in  std_logic;
    pdl13     : out std_logic;
    \-pdla5a\ : in  std_logic;
    \-pdla6a\ : in  std_logic;
    \-pdla7a\ : in  std_logic;
    \-pdla8a\ : in  std_logic;
    \-pdla9a\ : in  std_logic;
    \-pwpb\   : in  std_logic;
    l13       : in  std_logic;
    pdl12     : out std_logic;
    l12       : in  std_logic;
    pdl11     : out std_logic;
    l11       : in  std_logic;
    pdl10     : out std_logic;
    \-pwpc\   : in  std_logic;
    l10       : in  std_logic;
    pdl4      : out std_logic;
    l4        : in  std_logic;
    pdl3      : out std_logic;
    l3        : in  std_logic;
    pdl2      : out std_logic;
    l2        : in  std_logic;
    pdl1      : out std_logic;
    l1        : in  std_logic;
    pdl0      : out std_logic;
    l0        : in  std_logic;
    pdl15     : out std_logic;
    l15       : in  std_logic;
    pdl14     : out std_logic;
    l14       : in  std_logic;
    pdl9      : out std_logic;
    l9        : in  std_logic;
    pdl8      : out std_logic;
    l8        : in  std_logic;
    pdl7      : out std_logic;
    l7        : in  std_logic;
    pdl6      : out std_logic;
    l6        : in  std_logic;
    pdl5      : out std_logic;
    l5        : in  std_logic
    );
end;
