-- VMEM2 -- VIRTUAL MEMORY MAP STAGE 1

library work;
use work.dip.all;
use work.misc.all;

architecture behv of cadr_vmem2 is
begin
vmem2_1b01 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo20\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma20\);
vmem2_1b02 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo21\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma21\);
vmem2_1b03 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo22\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma22\);
vmem2_1b04 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo23\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma23\);
vmem2_1b06 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo16\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma16\);
vmem2_1b07 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo17\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma17\);
vmem2_1b08 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo18\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma18\);
vmem2_1b09 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo19\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma19\);
vmem2_1b11 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo12\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma12\);
vmem2_1b12 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo13\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma13\);
vmem2_1b13 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo14\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma14\);
vmem2_1b14 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => \-vmo15\, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => \-vma15\);
vmem2_1b17 : dip_93s48 port map (p1 => \-vmo17\, p2 => \-vmo18\, p3 => \-vmo19\, p4 => \-vmo20\, p5 => \-vmo21\, p6 => \-vmo22\, p7 => \-vmo23\, p9 => vmoparm, p10 => open, p11 => \-vmo12\, p12 => \-vmo13\, p13 => \-vmo14\, p14 => \-vmo15\, p15 => \-vmo16\);
vmem2_1c05 : dip_93425a port map (p1 => gnd, p2 => vmap4b, p3 => vmap3b, p4 => vmap2b, p5 => vmap1b, p6 => vmap0b, p7 => vmopar, p9 => \-mapi12b\, p10 => \-mapi11b\, p11 => \-mapi10b\, p12 => \-mapi9b\, p13 => \-mapi8b\, p14 => \-vm1wpb\, p15 => vm1pari);
vmem2_1c10 : dip_74s240 port map (p1 => gnd, p2 => '0', p3 => vmap0b, p4 => '0', p5 => vmap1b, p6 => '0', p7 => vmap2b, p8 => \-vmap4\, p9 => vmap3b, p11 => \-vmap3\, p12 => vmap4b, p13 => \-vmap2\, p14 => open, p15 => \-vmap1\, p16 => open, p17 => \-vmap0\, p18 => open, p19 => gnd);
vmem2_1d03 : dip_93s48 port map (p1 => \-vmo5\, p2 => \-vmo6\, p3 => \-vmo7\, p4 => \-vmo8\, p5 => \-vmo9\, p6 => \-vmo10\, p7 => \-vmo11\, p9 => vmoparl, p10 => open, p11 => \-vmo0\, p12 => \-vmo1\, p13 => \-vmo2\, p14 => \-vmo3\, p15 => \-vmo4\);
vmem2_1d12 : dip_74s86 port map (p1 => '0', p2 => '0', p3 => open, p4 => vmoparm, p5 => vmoparl, p6 => vmoparck, p8 => vmoparodd, p9 => vmopar, p10 => vmoparck, p11 => open, p12 => '0', p13 => '0');
end architecture;
