library ieee;
use ieee.std_logic_1164.all;

entity cadr_mskg4 is
  port (
    \a=m\   : inout std_logic;
    msk24   : inout std_logic;
    msk25   : inout std_logic;
    msk26   : inout std_logic;
    msk27   : inout std_logic;
    msk28   : inout std_logic;
    msk29   : inout std_logic;
    msk30   : inout std_logic;
    msk31   : inout std_logic;
    mskl0   : in  std_logic;
    mskl1   : in  std_logic;
    mskl2   : in  std_logic;
    mskl3   : in  std_logic;
    mskl4   : in  std_logic;
    gnd     : in  std_logic;
    mskr0   : in  std_logic;
    mskr1   : in  std_logic;
    mskr2   : in  std_logic;
    mskr3   : in  std_logic;
    mskr4   : in  std_logic;
    msk8    : inout std_logic;
    msk9    : inout std_logic;
    msk10   : inout std_logic;
    msk11   : inout std_logic;
    msk12   : inout std_logic;
    msk13   : inout std_logic;
    msk14   : inout std_logic;
    msk15   : inout std_logic;
    ir31    : in  std_logic;
    \-ir31\ : out std_logic;
    ir13    : in  std_logic;
    \-ir13\ : out std_logic;
    \-ir12\ : out std_logic;
    ir12    : in  std_logic;
    msk16   : inout std_logic;
    msk17   : inout std_logic;
    msk18   : inout std_logic;
    msk19   : inout std_logic;
    msk20   : inout std_logic;
    msk21   : inout std_logic;
    msk22   : inout std_logic;
    msk23   : inout std_logic;
    aeqm    : out std_logic;
    msk0    : inout std_logic;
    msk1    : inout std_logic;
    msk2    : inout std_logic;
    msk3    : inout std_logic;
    msk4    : inout std_logic;
    msk5    : inout std_logic;
    msk6    : inout std_logic;
    msk7    : inout std_logic);
end;
