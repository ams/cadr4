library ieee;
use ieee.std_logic_1164.all;

entity cadr_ior is
  port (
    i12   : in  std_logic;
    ob12  : in  std_logic;
    iob12 : out std_logic;
    i13   : in  std_logic;
    ob13  : in  std_logic;
    iob13 : out std_logic;
    iob14 : out std_logic;
    i14   : in  std_logic;
    ob14  : in  std_logic;
    iob15 : out std_logic;
    i15   : in  std_logic;
    ob15  : in  std_logic;
    i8    : in  std_logic;
    ob8   : in  std_logic;
    iob8  : out std_logic;
    i9    : in  std_logic;
    ob9   : in  std_logic;
    iob9  : out std_logic;
    iob10 : out std_logic;
    i10   : in  std_logic;
    ob10  : in  std_logic;
    iob11 : out std_logic;
    i11   : in  std_logic;
    ob11  : in  std_logic;
    i4    : in  std_logic;
    ob4   : in  std_logic;
    iob4  : out std_logic;
    i5    : in  std_logic;
    ob5   : in  std_logic;
    iob5  : out std_logic;
    iob6  : out std_logic;
    i6    : in  std_logic;
    ob6   : in  std_logic;
    iob7  : out std_logic;
    i7    : in  std_logic;
    ob7   : in  std_logic;
    i0    : in  std_logic;
    ob0   : in  std_logic;
    iob0  : out std_logic;
    i1    : in  std_logic;
    ob1   : in  std_logic;
    iob1  : out std_logic;
    iob2  : out std_logic;
    i2    : in  std_logic;
    ob2   : in  std_logic;
    iob3  : out std_logic;
    i3    : in  std_logic;
    ob3   : in  std_logic;
    i20   : in  std_logic;
    ob20  : in  std_logic;
    iob20 : out std_logic;
    i21   : in  std_logic;
    ob21  : in  std_logic;
    iob21 : out std_logic;
    iob22 : out std_logic;
    i22   : in  std_logic;
    ob22  : in  std_logic;
    iob23 : out std_logic;
    i23   : in  std_logic;
    ob23  : in  std_logic;
    i16   : in  std_logic;
    ob16  : in  std_logic;
    iob16 : out std_logic;
    i17   : in  std_logic;
    ob17  : in  std_logic;
    iob17 : out std_logic;
    iob18 : out std_logic;
    i18   : in  std_logic;
    ob18  : in  std_logic;
    iob19 : out std_logic;
    i19   : in  std_logic;
    ob19  : in  std_logic;
    i44   : in  std_logic;
    iob44 : out std_logic;
    i45   : in  std_logic;
    iob45 : out std_logic;
    iob46 : out std_logic;
    i46   : in  std_logic;
    iob47 : out std_logic;
    i47   : in  std_logic;
    i40   : in  std_logic;
    iob40 : out std_logic;
    i41   : in  std_logic;
    iob41 : out std_logic;
    iob42 : out std_logic;
    i42   : in  std_logic;
    iob43 : out std_logic;
    i43   : in  std_logic;
    i36   : in  std_logic;
    iob36 : out std_logic;
    i37   : in  std_logic;
    iob37 : out std_logic;
    iob38 : out std_logic;
    i38   : in  std_logic;
    iob39 : out std_logic;
    i39   : in  std_logic;
    i32   : in  std_logic;
    iob32 : out std_logic;
    i33   : in  std_logic;
    iob33 : out std_logic;
    iob34 : out std_logic;
    i34   : in  std_logic;
    iob35 : out std_logic;
    i35   : in  std_logic;
    i28   : in  std_logic;
    iob28 : out std_logic;
    i29   : in  std_logic;
    iob29 : out std_logic;
    iob30 : out std_logic;
    i30   : in  std_logic;
    iob31 : out std_logic;
    i31   : in  std_logic;
    i24   : in  std_logic;
    ob24  : in  std_logic;
    iob24 : out std_logic;
    i25   : in  std_logic;
    ob25  : in  std_logic;
    iob25 : out std_logic;
    iob26 : out std_logic;
    i26   : in  std_logic;
    iob27 : out std_logic;
    i27   : in  std_logic);
end;
