library ieee;
use ieee.std_logic_1164.all;

entity busint_uba is
  port (
    \-ubadrive\     : in     std_logic;
    \c1 out\        : in     std_logic;
    uao1            : in     std_logic;
    uao10           : in     std_logic;
    uao11           : in     std_logic;
    uao12           : in     std_logic;
    uao13           : in     std_logic;
    uao14           : in     std_logic;
    uao15           : in     std_logic;
    uao16           : in     std_logic;
    uao17           : in     std_logic;
    uao2            : in     std_logic;
    uao3            : in     std_logic;
    uao4            : in     std_logic;
    uao5            : in     std_logic;
    uao6            : in     std_logic;
    uao7            : in     std_logic;
    uao8            : in     std_logic;
    uao9            : in     std_logic;
    \-ub adr0\      : inout  std_logic;
    \-ub adr10\     : inout  std_logic;
    \-ub adr11\     : inout  std_logic;
    \-ub adr12\     : inout  std_logic;
    \-ub adr13\     : inout  std_logic;
    \-ub adr14\     : inout  std_logic;
    \-ub adr15\     : inout  std_logic;
    \-ub adr16\     : inout  std_logic;
    \-ub adr17\     : inout  std_logic;
    \-ub adr1\      : inout  std_logic;
    \-ub adr2\      : inout  std_logic;
    \-ub adr3\      : inout  std_logic;
    \-ub adr4\      : inout  std_logic;
    \-ub adr5\      : inout  std_logic;
    \-ub adr6\      : inout  std_logic;
    \-ub adr7\      : inout  std_logic;
    \-ub adr8\      : inout  std_logic;
    \-ub adr9\      : inout  std_logic;
    \-ub c1\        : inout  std_logic;
    \-uba 12\       : out    std_logic;
    \-uba 14\       : out    std_logic;
    \-uba 15\       : out    std_logic;
    \-uba 7\        : out    std_logic;
    \-uba 8\        : out    std_logic;
    \-uba 9\        : out    std_logic;
    \c1 in\         : out    std_logic;
    uba0            : out    std_logic;
    uba1            : out    std_logic;
    uba10           : out    std_logic;
    uba11           : out    std_logic;
    uba12           : out    std_logic;
    uba13           : out    std_logic;
    uba14           : out    std_logic;
    uba15           : out    std_logic;
    uba16           : out    std_logic;
    uba17           : out    std_logic;
    uba2            : out    std_logic;
    uba3            : out    std_logic;
    uba4            : out    std_logic;
    uba5            : out    std_logic;
    uba6            : out    std_logic;
    uba7            : out    std_logic;
    uba8            : out    std_logic;
    uba9            : out    std_logic
  );
end entity;
