library ieee;
use ieee.std_logic_1164.all;

entity cadr_shift0 is
  port (
    \-s4\           : in     std_logic;
    m0              : in     std_logic;
    m1              : in     std_logic;
    m10             : in     std_logic;
    m11             : in     std_logic;
    m12             : in     std_logic;
    m13             : in     std_logic;
    m14             : in     std_logic;
    m15             : in     std_logic;
    m2              : in     std_logic;
    m29             : in     std_logic;
    m3              : in     std_logic;
    m30             : in     std_logic;
    m31             : in     std_logic;
    m4              : in     std_logic;
    m5              : in     std_logic;
    m6              : in     std_logic;
    m7              : in     std_logic;
    m8              : in     std_logic;
    m9              : in     std_logic;
    s0              : in     std_logic;
    s1              : in     std_logic;
    s2a             : in     std_logic;
    s3a             : in     std_logic;
    s4              : in     std_logic;
    sa16            : in     std_logic;
    sa17            : in     std_logic;
    sa18            : in     std_logic;
    sa19            : in     std_logic;
    sa20            : in     std_logic;
    sa21            : in     std_logic;
    sa22            : in     std_logic;
    sa23            : in     std_logic;
    sa24            : in     std_logic;
    sa25            : in     std_logic;
    sa26            : in     std_logic;
    sa27            : in     std_logic;
    sa28            : in     std_logic;
    sa29            : in     std_logic;
    sa30            : in     std_logic;
    sa31            : in     std_logic;
    r0              : out    std_logic;
    r1              : out    std_logic;
    r10             : out    std_logic;
    r11             : out    std_logic;
    r12             : out    std_logic;
    r13             : out    std_logic;
    r14             : out    std_logic;
    r15             : out    std_logic;
    r2              : out    std_logic;
    r3              : out    std_logic;
    r4              : out    std_logic;
    r5              : out    std_logic;
    r6              : out    std_logic;
    r7              : out    std_logic;
    r8              : out    std_logic;
    r9              : out    std_logic;
    sa0             : out    std_logic;
    sa1             : out    std_logic;
    sa10            : out    std_logic;
    sa11            : out    std_logic;
    sa12            : out    std_logic;
    sa13            : out    std_logic;
    sa14            : out    std_logic;
    sa15            : out    std_logic;
    sa2             : out    std_logic;
    sa3             : out    std_logic;
    sa4             : out    std_logic;
    sa5             : out    std_logic;
    sa6             : out    std_logic;
    sa7             : out    std_logic;
    sa8             : out    std_logic;
    sa9             : out    std_logic
  );
end entity cadr_shift0;
