library ieee;
use ieee.std_logic_1164.all;

entity busint_ubxa is
  port (
    \-ubaddr>xbus\  : in     std_logic;
    uba2            : in     std_logic;
    uba3            : in     std_logic;
    uba4            : in     std_logic;
    uba5            : in     std_logic;
    uba6            : in     std_logic;
    uba7            : in     std_logic;
    uba8            : in     std_logic;
    uba9            : in     std_logic;
    ubma10          : in     std_logic;
    ubma11          : in     std_logic;
    ubma12          : in     std_logic;
    ubma13          : in     std_logic;
    ubma14          : in     std_logic;
    ubma15          : in     std_logic;
    ubma16          : in     std_logic;
    ubma17          : in     std_logic;
    ubma18          : in     std_logic;
    ubma19          : in     std_logic;
    ubma20          : in     std_logic;
    ubma21          : in     std_logic;
    ubma8           : in     std_logic;
    ubma9           : in     std_logic;
    xao0            : out    std_logic;
    xao1            : out    std_logic;
    xao10           : out    std_logic;
    xao11           : out    std_logic;
    xao12           : out    std_logic;
    xao13           : out    std_logic;
    xao14           : out    std_logic;
    xao15           : out    std_logic;
    xao16           : out    std_logic;
    xao17           : out    std_logic;
    xao18           : out    std_logic;
    xao19           : out    std_logic;
    xao2            : out    std_logic;
    xao20           : out    std_logic;
    xao21           : out    std_logic;
    xao3            : out    std_logic;
    xao4            : out    std_logic;
    xao5            : out    std_logic;
    xao6            : out    std_logic;
    xao7            : out    std_logic;
    xao8            : out    std_logic;
    xao9            : out    std_logic
  );
end entity busint_ubxa;
