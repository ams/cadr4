library ieee;
use ieee.std_logic_1164.all;

entity cadr_vmem1 is
  port (
    \-vm1wpa\       : in     std_logic;
    \-vma0\         : in     std_logic;
    \-vma10\        : in     std_logic;
    \-vma11\        : in     std_logic;
    \-vma12\        : in     std_logic;
    \-vma13\        : in     std_logic;
    \-vma14\        : in     std_logic;
    \-vma15\        : in     std_logic;
    \-vma16\        : in     std_logic;
    \-vma17\        : in     std_logic;
    \-vma18\        : in     std_logic;
    \-vma19\        : in     std_logic;
    \-vma1\         : in     std_logic;
    \-vma20\        : in     std_logic;
    \-vma21\        : in     std_logic;
    \-vma22\        : in     std_logic;
    \-vma23\        : in     std_logic;
    \-vma2\         : in     std_logic;
    \-vma3\         : in     std_logic;
    \-vma4\         : in     std_logic;
    \-vma5\         : in     std_logic;
    \-vma6\         : in     std_logic;
    \-vma7\         : in     std_logic;
    \-vma8\         : in     std_logic;
    \-vma9\         : in     std_logic;
    \-vmap0\        : in     std_logic;
    \-vmap1\        : in     std_logic;
    \-vmap2\        : in     std_logic;
    \-vmap3\        : in     std_logic;
    \-vmap4\        : in     std_logic;
    mapi10          : in     std_logic;
    mapi11          : in     std_logic;
    mapi12          : in     std_logic;
    mapi8           : in     std_logic;
    mapi9           : in     std_logic;
    \-mapi10a\      : out    std_logic;
    \-mapi10b\      : out    std_logic;
    \-mapi11a\      : out    std_logic;
    \-mapi11b\      : out    std_logic;
    \-mapi12a\      : out    std_logic;
    \-mapi12b\      : out    std_logic;
    \-mapi8a\       : out    std_logic;
    \-mapi8b\       : out    std_logic;
    \-mapi9a\       : out    std_logic;
    \-mapi9b\       : out    std_logic;
    \-vm1lpar\      : out    std_logic;
    \-vmo0\         : out    std_logic;
    \-vmo10\        : out    std_logic;
    \-vmo11\        : out    std_logic;
    \-vmo1\         : out    std_logic;
    \-vmo2\         : out    std_logic;
    \-vmo3\         : out    std_logic;
    \-vmo4\         : out    std_logic;
    \-vmo5\         : out    std_logic;
    \-vmo6\         : out    std_logic;
    \-vmo7\         : out    std_logic;
    \-vmo8\         : out    std_logic;
    \-vmo9\         : out    std_logic;
    vm1mpar         : out    std_logic;
    vm1pari         : out    std_logic;
    vmap0a          : out    std_logic;
    vmap1a          : out    std_logic;
    vmap2a          : out    std_logic;
    vmap3a          : out    std_logic;
    vmap4a          : out    std_logic
  );
end entity cadr_vmem1;
