library ieee;
use ieee.std_logic_1164.all;

entity cadr_spcw is
  port (
    destspcd : in  std_logic;
    reta12   : out std_logic;
    l12      : in  std_logic;
    spcw12   : out std_logic;
    reta13   : out std_logic;
    l13      : in  std_logic;
    spcw13   : out std_logic;
    spcw14   : out std_logic;
    l14      : in  std_logic;
    gnd      : in  std_logic;
    spcw15   : out std_logic;
    l15      : in  std_logic;
    reta8    : out std_logic;
    l8       : in  std_logic;
    spcw8    : out std_logic;
    reta9    : out std_logic;
    l9       : in  std_logic;
    spcw9    : out std_logic;
    spcw10   : out std_logic;
    l10      : in  std_logic;
    reta10   : out std_logic;
    spcw11   : out std_logic;
    l11      : in  std_logic;
    reta11   : out std_logic;
    reta4    : out std_logic;
    l4       : in  std_logic;
    spcw4    : out std_logic;
    reta5    : out std_logic;
    l5       : in  std_logic;
    spcw5    : out std_logic;
    spcw6    : out std_logic;
    l6       : in  std_logic;
    reta6    : out std_logic;
    spcw7    : out std_logic;
    l7       : in  std_logic;
    reta7    : out std_logic;
    reta0    : out std_logic;
    l0       : in  std_logic;
    spcw0    : out std_logic;
    reta1    : out std_logic;
    l1       : in  std_logic;
    spcw1    : out std_logic;
    spcw2    : out std_logic;
    l2       : in  std_logic;
    reta2    : out std_logic;
    spcw3    : out std_logic;
    l3       : in  std_logic;
    reta3    : out std_logic;
    n        : in  std_logic;
    ipc12    : in  std_logic;
    wpc12    : in  std_logic;
    wpc13    : in  std_logic;
    ipc13    : in  std_logic;
    clk4d    : in  std_logic;
    ipc8     : in  std_logic;
    wpc8     : in  std_logic;
    wpc9     : in  std_logic;
    ipc9     : in  std_logic;
    ipc10    : in  std_logic;
    wpc10    : in  std_logic;
    wpc11    : in  std_logic;
    ipc11    : in  std_logic;
    ipc4     : in  std_logic;
    wpc4     : in  std_logic;
    wpc5     : in  std_logic;
    ipc5     : in  std_logic;
    ipc6     : in  std_logic;
    wpc6     : in  std_logic;
    wpc7     : in  std_logic;
    ipc7     : in  std_logic;
    ipc0     : in  std_logic;
    wpc0     : in  std_logic;
    wpc1     : in  std_logic;
    ipc1     : in  std_logic;
    ipc2     : in  std_logic;
    wpc2     : in  std_logic;
    wpc3     : in  std_logic;
    ipc3     : in  std_logic;
    l16      : in  std_logic;
    spcw16   : out std_logic;
    l17      : in  std_logic;
    spcw17   : out std_logic;
    spcw18   : out std_logic;
    l18      : in  std_logic
    );
end;
