library ieee;
use ieee.std_logic_1164.all;

entity cadr_iwr is
  port (
    gnd   : in  std_logic;
    iwr47 : out std_logic;
    aa15  : in  std_logic;
    aa14  : in  std_logic;
    iwr46 : out std_logic;
    iwr45 : out std_logic;
    aa13  : in  std_logic;
    aa12  : in  std_logic;
    iwr44 : out std_logic;
    clk2c : in  std_logic;
    iwr43 : out std_logic;
    aa11  : in  std_logic;
    aa10  : in  std_logic;
    iwr42 : out std_logic;
    iwr41 : out std_logic;
    aa9   : in  std_logic;
    aa8   : in  std_logic;
    iwr40 : out std_logic;
    iwr39 : out std_logic;
    aa7   : in  std_logic;
    aa6   : in  std_logic;
    iwr38 : out std_logic;
    iwr37 : out std_logic;
    aa5   : in  std_logic;
    aa4   : in  std_logic;
    iwr36 : out std_logic;
    iwr35 : out std_logic;
    aa3   : in  std_logic;
    aa2   : in  std_logic;
    iwr34 : out std_logic;
    iwr33 : out std_logic;
    aa1   : in  std_logic;
    aa0   : in  std_logic;
    iwr32 : out std_logic;
    iwr15 : out std_logic;
    m15   : in  std_logic;
    m14   : in  std_logic;
    iwr14 : out std_logic;
    iwr13 : out std_logic;
    m13   : in  std_logic;
    m12   : in  std_logic;
    iwr12 : out std_logic;
    clk4c : in  std_logic;
    iwr11 : out std_logic;
    m11   : in  std_logic;
    m10   : in  std_logic;
    iwr10 : out std_logic;
    iwr9  : out std_logic;
    m9    : in  std_logic;
    m8    : in  std_logic;
    iwr8  : out std_logic;
    iwr7  : out std_logic;
    m7    : in  std_logic;
    m6    : in  std_logic;
    iwr6  : out std_logic;
    iwr5  : out std_logic;
    m5    : in  std_logic;
    m4    : in  std_logic;
    iwr4  : out std_logic;
    iwr3  : out std_logic;
    m3    : in  std_logic;
    m2    : in  std_logic;
    iwr2  : out std_logic;
    iwr1  : out std_logic;
    m1    : in  std_logic;
    m0    : in  std_logic;
    iwr0  : out std_logic;
    iwr31 : out std_logic;
    m31   : in  std_logic;
    m30   : in  std_logic;
    iwr30 : out std_logic;
    iwr29 : out std_logic;
    m29   : in  std_logic;
    m28   : in  std_logic;
    iwr28 : out std_logic;
    iwr27 : out std_logic;
    m27   : in  std_logic;
    m26   : in  std_logic;
    iwr26 : out std_logic;
    iwr25 : out std_logic;
    m25   : in  std_logic;
    m24   : in  std_logic;
    iwr24 : out std_logic;
    iwr23 : out std_logic;
    m23   : in  std_logic;
    m22   : in  std_logic;
    iwr22 : out std_logic;
    iwr21 : out std_logic;
    m21   : in  std_logic;
    m20   : in  std_logic;
    iwr20 : out std_logic;
    iwr19 : out std_logic;
    m19   : in  std_logic;
    m18   : in  std_logic;
    iwr18 : out std_logic;
    iwr17 : out std_logic;
    m17   : in  std_logic;
    m16   : in  std_logic;
    iwr16 : out std_logic
    );
end;
