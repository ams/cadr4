library ieee;
use ieee.std_logic_1164.all;

entity cadr_spy2 is
  port (
    \-spy.al\    : out std_logic;
    aa15         : in  std_logic;
    spy8         : out std_logic;
    aa14         : in  std_logic;
    spy9         : out std_logic;
    aa13         : in  std_logic;
    spy10        : out std_logic;
    aa12         : in  std_logic;
    spy11        : out std_logic;
    aa11         : in  std_logic;
    spy12        : out std_logic;
    aa10         : in  std_logic;
    spy13        : out std_logic;
    aa9          : in  std_logic;
    spy14        : out std_logic;
    aa8          : in  std_logic;
    spy15        : out std_logic;
    aa7          : in  std_logic;
    spy0         : out std_logic;
    aa6          : in  std_logic;
    spy1         : out std_logic;
    aa5          : in  std_logic;
    spy2         : out std_logic;
    aa4          : in  std_logic;
    spy3         : out std_logic;
    aa3          : in  std_logic;
    spy4         : out std_logic;
    aa2          : in  std_logic;
    spy5         : out std_logic;
    aa1          : in  std_logic;
    spy6         : out std_logic;
    aa0          : in  std_logic;
    spy7         : out std_logic;
    \-spy.ah\    : in  std_logic;
    a31a         : in  std_logic;
    a30          : in  std_logic;
    a29          : in  std_logic;
    a28          : in  std_logic;
    a27          : in  std_logic;
    a26          : in  std_logic;
    a25          : in  std_logic;
    a24          : in  std_logic;
    a23          : in  std_logic;
    a22          : in  std_logic;
    a21          : in  std_logic;
    a20          : in  std_logic;
    a19          : in  std_logic;
    a18          : in  std_logic;
    a17          : in  std_logic;
    a16          : in  std_logic;
    \-spy.flag2\ : in  std_logic;
    ir48         : in  std_logic;
    nop          : in  std_logic;
    \-vmaok\     : in  std_logic;
    jcond        : in  std_logic;
    pcs1         : in  std_logic;
    pcs0         : in  std_logic;
    wmapd        : in  std_logic;
    destspcd     : in  std_logic;
    iwrited      : in  std_logic;
    imodd        : in  std_logic;
    pdlwrited    : in  std_logic;
    spushd       : in  std_logic;
    \-spy.ml\    : in  std_logic;
    m15          : in  std_logic;
    m14          : in  std_logic;
    m13          : in  std_logic;
    m12          : in  std_logic;
    m11          : in  std_logic;
    m10          : in  std_logic;
    m9           : in  std_logic;
    m8           : in  std_logic;
    m7           : in  std_logic;
    m6           : in  std_logic;
    m5           : in  std_logic;
    m4           : in  std_logic;
    m3           : in  std_logic;
    m2           : in  std_logic;
    m1           : in  std_logic;
    m0           : in  std_logic;
    \-spy.mh\    : in  std_logic;
    m23          : in  std_logic;
    m22          : in  std_logic;
    m21          : in  std_logic;
    m20          : in  std_logic;
    m19          : in  std_logic;
    m18          : in  std_logic;
    m17          : in  std_logic;
    m16          : in  std_logic;
    m31          : in  std_logic;
    m30          : in  std_logic;
    m29          : in  std_logic;
    m28          : in  std_logic;
    m27          : in  std_logic;
    m26          : in  std_logic;
    m25          : in  std_logic;
    m24          : in  std_logic);
end;
