library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_7420 is
  port (
    g1a   : in  std_logic;
    g1b   : in  std_logic;
    g1c   : in  std_logic;
    g1d   : in  std_logic;
    g1y_n : out std_logic;
    g2y_n : out std_logic;
    g2a   : in  std_logic;
    g2b   : in  std_logic;
    g2c   : in  std_logic;
    g2d   : in  std_logic
    );
end ic_7420;

architecture ttl of ic_7420 is
begin

end ttl;
