library ieee;
use ieee.std_logic_1164.all;

entity cadr_trap is
  port (
    \-md0\          : in     std_logic;
    \-md10\         : in     std_logic;
    \-md11\         : in     std_logic;
    \-md12\         : in     std_logic;
    \-md13\         : in     std_logic;
    \-md14\         : in     std_logic;
    \-md15\         : in     std_logic;
    \-md16\         : in     std_logic;
    \-md17\         : in     std_logic;
    \-md18\         : in     std_logic;
    \-md19\         : in     std_logic;
    \-md1\          : in     std_logic;
    \-md20\         : in     std_logic;
    \-md21\         : in     std_logic;
    \-md22\         : in     std_logic;
    \-md23\         : in     std_logic;
    \-md24\         : in     std_logic;
    \-md25\         : in     std_logic;
    \-md26\         : in     std_logic;
    \-md27\         : in     std_logic;
    \-md28\         : in     std_logic;
    \-md29\         : in     std_logic;
    \-md2\          : in     std_logic;
    \-md30\         : in     std_logic;
    \-md31\         : in     std_logic;
    \-md3\          : in     std_logic;
    \-md4\          : in     std_logic;
    \-md5\          : in     std_logic;
    \-md6\          : in     std_logic;
    \-md7\          : in     std_logic;
    \-md8\          : in     std_logic;
    \-md9\          : in     std_logic;
    \-wait\         : in     std_logic;
    \boot.trap\     : in     std_logic;
    \use.md\        : in     std_logic;
    mdhaspar        : in     std_logic;
    mdpar           : in     std_logic;
    trapenb         : in     std_logic;
    \-memparok\     : out    std_logic;
    \-parerr\       : out    std_logic;
    \-trap\         : out    std_logic;
    \-trapenb\      : out    std_logic;
    mdparerr        : out    std_logic;
    mdpareven       : out    std_logic;
    mdparl          : out    std_logic;
    mdparm          : out    std_logic;
    mdparodd        : out    std_logic;
    memparok        : out    std_logic;
    trapa           : out    std_logic;
    trapb           : out    std_logic
  );
end entity cadr_trap;
