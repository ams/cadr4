library ieee;
use ieee.std_logic_1164.all;

entity alu1 is
  port (
    a31a     : in  std_logic;
    m31b     : out std_logic;
    aluf3a   : in  std_logic;
    aluf2a   : in  std_logic;
    aluf1a   : in  std_logic;
    aluf0a   : in  std_logic;
    \-cin32\ : in  std_logic;
    alumode  : in  std_logic;
    alu32    : out std_logic;
    m31      : in  std_logic;
    hi12     : in  std_logic;
    a28      : in  std_logic;
    m28      : in  std_logic;
    \-cin28\ : in  std_logic;
    alu28    : out std_logic;
    alu29    : out std_logic;
    alu30    : out std_logic;
    alu31    : out std_logic;
    aeqm     : out std_logic;
    xout31   : out std_logic;
    yout31   : out std_logic;
    a31b     : in  std_logic;
    a30      : in  std_logic;
    m30      : in  std_logic;
    a29      : in  std_logic;
    m29      : in  std_logic;
    a20      : in  std_logic;
    m20      : in  std_logic;
    \-cin20\ : in  std_logic;
    alu20    : out std_logic;
    alu21    : out std_logic;
    alu22    : out std_logic;
    alu23    : out std_logic;
    xout23   : out std_logic;
    yout23   : out std_logic;
    a23      : in  std_logic;
    m23      : in  std_logic;
    a22      : in  std_logic;
    m22      : in  std_logic;
    a21      : in  std_logic;
    m21      : in  std_logic;
    a24      : in  std_logic;
    m24      : in  std_logic;
    \-cin24\ : in  std_logic;
    alu24    : out std_logic;
    alu25    : out std_logic;
    alu26    : out std_logic;
    alu27    : out std_logic;
    xout27   : out std_logic;
    yout27   : out std_logic;
    a27      : in  std_logic;
    m27      : in  std_logic;
    a26      : in  std_logic;
    m26      : in  std_logic;
    a25      : in  std_logic;
    m25      : in  std_logic;
    a16      : in  std_logic;
    m16      : in  std_logic;
    \-cin16\ : in  std_logic;
    alu16    : out std_logic;
    alu17    : out std_logic;
    alu18    : out std_logic;
    alu19    : out std_logic;
    xout19   : out std_logic;
    yout19   : out std_logic;
    a19      : in  std_logic;
    m19      : in  std_logic;
    a18      : in  std_logic;
    m18      : in  std_logic;
    a17      : in  std_logic;
    m17      : in  std_logic);
end;
