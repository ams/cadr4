library ieee;
use ieee.std_logic_1164.all;

entity cadr_q is
  port (
    hi7      : in  std_logic;
    q23      : out std_logic;
    alu24    : in  std_logic;
    alu25    : in  std_logic;
    alu26    : in  std_logic;
    alu27    : in  std_logic;
    q28      : out std_logic;
    qs0      : in  std_logic;
    qs1      : in  std_logic;
    clk2b    : in  std_logic;
    q27      : out std_logic;
    q26      : out std_logic;
    q25      : out std_logic;
    q24      : out std_logic;
    alu28    : in  std_logic;
    alu29    : in  std_logic;
    alu30    : in  std_logic;
    alu31    : in  std_logic;
    alu0     : in  std_logic;
    q31      : out std_logic;
    q30      : out std_logic;
    q29      : out std_logic;
    q15      : out std_logic;
    alu16    : in  std_logic;
    alu17    : in  std_logic;
    alu18    : in  std_logic;
    alu19    : in  std_logic;
    q20      : out std_logic;
    q19      : out std_logic;
    q18      : out std_logic;
    q17      : out std_logic;
    q16      : out std_logic;
    alu20    : in  std_logic;
    alu21    : in  std_logic;
    alu22    : in  std_logic;
    alu23    : in  std_logic;
    q22      : out std_logic;
    q21      : out std_logic;
    q7       : out std_logic;
    alu8     : in  std_logic;
    alu9     : in  std_logic;
    alu10    : in  std_logic;
    alu11    : in  std_logic;
    q12      : out std_logic;
    q11      : out std_logic;
    q10      : out std_logic;
    q9       : out std_logic;
    q8       : out std_logic;
    alu12    : in  std_logic;
    alu13    : in  std_logic;
    alu14    : in  std_logic;
    alu15    : in  std_logic;
    q14      : out std_logic;
    q13      : out std_logic;
    \-alu31\ : in  std_logic;
    alu1     : in  std_logic;
    alu2     : in  std_logic;
    alu3     : in  std_logic;
    q4       : out std_logic;
    q3       : out std_logic;
    q2       : out std_logic;
    q1       : out std_logic;
    q0       : out std_logic;
    alu4     : in  std_logic;
    alu5     : in  std_logic;
    alu6     : in  std_logic;
    alu7     : in  std_logic;
    q6       : out std_logic;
    q5       : out std_logic);
end;
