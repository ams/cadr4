library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_ireg is
  port (
    \-destimod0\ : in  std_logic;
    ir15         : out std_logic;
    iob15        : in  std_logic;
    i15          : in  std_logic;
    i14          : in  std_logic;
    iob14        : in  std_logic;
    ir14         : out std_logic;
    clk3a        : in  std_logic;
    ir13         : out std_logic;
    iob13        : in  std_logic;
    i13          : in  std_logic;
    i12          : in  std_logic;
    iob12        : in  std_logic;
    ir12         : out std_logic;
    ir11         : out std_logic;
    iob11        : in  std_logic;
    i11          : in  std_logic;
    i10          : in  std_logic;
    iob10        : in  std_logic;
    ir10         : out std_logic;
    ir9          : out std_logic;
    iob9         : in  std_logic;
    i9           : in  std_logic;
    i8           : in  std_logic;
    iob8         : in  std_logic;
    ir8          : out std_logic;
    ir7          : out std_logic;
    iob7         : in  std_logic;
    i7           : in  std_logic;
    i6           : in  std_logic;
    iob6         : in  std_logic;
    ir6          : out std_logic;
    ir5          : out std_logic;
    iob5         : in  std_logic;
    i5           : in  std_logic;
    i4           : in  std_logic;
    iob4         : in  std_logic;
    ir4          : out std_logic;
    ir3          : out std_logic;
    iob3         : in  std_logic;
    i3           : in  std_logic;
    i2           : in  std_logic;
    iob2         : in  std_logic;
    ir2          : out std_logic;
    ir1          : out std_logic;
    iob1         : in  std_logic;
    i1           : in  std_logic;
    i0           : in  std_logic;
    iob0         : in  std_logic;
    ir0          : out std_logic;
    ir23         : out std_logic;
    iob23        : in  std_logic;
    i23          : in  std_logic;
    i22          : in  std_logic;
    iob22        : in  std_logic;
    ir22         : out std_logic;
    clk3b        : in  std_logic;
    ir21         : out std_logic;
    iob21        : in  std_logic;
    i21          : in  std_logic;
    i20          : in  std_logic;
    iob20        : in  std_logic;
    ir20         : out std_logic;
    ir19         : out std_logic;
    iob19        : in  std_logic;
    i19          : in  std_logic;
    i18          : in  std_logic;
    iob18        : in  std_logic;
    ir18         : out std_logic;
    ir17         : out std_logic;
    iob17        : in  std_logic;
    i17          : in  std_logic;
    i16          : in  std_logic;
    iob16        : in  std_logic;
    ir16         : out std_logic;
    \-destimod1\ : in  std_logic;
    i48          : in  std_logic;
    gnd          : in  std_logic;
    ir48         : out std_logic;
    ir47         : out std_logic;
    iob47        : in  std_logic;
    i47          : in  std_logic;
    i46          : in  std_logic;
    iob46        : in  std_logic;
    ir46         : out std_logic;
    ir45         : out std_logic;
    iob45        : in  std_logic;
    i45          : in  std_logic;
    i44          : in  std_logic;
    iob44        : in  std_logic;
    ir44         : out std_logic;
    ir43         : out std_logic;
    iob43        : in  std_logic;
    i43          : in  std_logic;
    i42          : in  std_logic;
    iob42        : in  std_logic;
    ir42         : out std_logic;
    ir41         : out std_logic;
    iob41        : in  std_logic;
    i41          : in  std_logic;
    i40          : in  std_logic;
    iob40        : in  std_logic;
    ir40         : out std_logic;
    ir39         : out std_logic;
    iob39        : in  std_logic;
    i39          : in  std_logic;
    i38          : in  std_logic;
    iob38        : in  std_logic;
    ir38         : out std_logic;
    ir37         : out std_logic;
    iob37        : in  std_logic;
    i37          : in  std_logic;
    i36          : in  std_logic;
    iob36        : in  std_logic;
    ir36         : out std_logic;
    ir35         : out std_logic;
    iob35        : in  std_logic;
    i35          : in  std_logic;
    i34          : in  std_logic;
    iob34        : in  std_logic;
    ir34         : out std_logic;
    ir33         : out std_logic;
    iob33        : in  std_logic;
    i33          : in  std_logic;
    i32          : in  std_logic;
    iob32        : in  std_logic;
    ir32         : out std_logic;
    ir31         : out std_logic;
    iob31        : in  std_logic;
    i31          : in  std_logic;
    i30          : in  std_logic;
    iob30        : in  std_logic;
    ir30         : out std_logic;
    ir29         : out std_logic;
    iob29        : in  std_logic;
    i29          : in  std_logic;
    i28          : in  std_logic;
    iob28        : in  std_logic;
    ir28         : out std_logic;
    ir27         : out std_logic;
    iob27        : in  std_logic;
    i27          : in  std_logic;
    i26          : in  std_logic;
    iob26        : in  std_logic;
    ir26         : out std_logic;
    ir25         : out std_logic;
    iob25        : in  std_logic;
    i25          : in  std_logic;
    i24          : in  std_logic;
    iob24        : in  std_logic;
    ir24         : out std_logic);
end;

architecture ttl of cadr4_ireg is
  signal nc371 : std_logic;
  signal nc372 : std_logic;
  signal nc373 : std_logic;
  signal nc374 : std_logic;
  signal nc375 : std_logic;
  signal nc376 : std_logic;
  signal nc377 : std_logic;
  signal nc378 : std_logic;
  signal nc379 : std_logic;
begin
  ireg_3c01 : am25s09 port map(sel => \-destimod0\, aq => ir15, a0 => iob15, a1 => i15, b1 => i14, b0 => iob14, bq => ir14, clk => clk3a, cq => ir13, c0 => iob13, c1 => i13, d1 => i12, d0 => iob12, dq => ir12);
  ireg_3c02 : am25s09 port map(sel => \-destimod0\, aq => ir11, a0 => iob11, a1 => i11, b1 => i10, b0 => iob10, bq => ir10, clk => clk3a, cq => ir9, c0 => iob9, c1 => i9, d1 => i8, d0 => iob8, dq => ir8);
  ireg_3c03 : am25s09 port map(sel => \-destimod0\, aq => ir7, a0 => iob7, a1 => i7, b1 => i6, b0 => iob6, bq => ir6, clk => clk3a, cq => ir5, c0 => iob5, c1 => i5, d1 => i4, d0 => iob4, dq => ir4);
  ireg_3c04 : am25s09 port map(sel => \-destimod0\, aq => ir3, a0 => iob3, a1 => i3, b1 => i2, b0 => iob2, bq => ir2, clk => clk3a, cq => ir1, c0 => iob1, c1 => i1, d1 => i0, d0 => iob0, dq => ir0);
  ireg_3c17 : am25s09 port map(sel => \-destimod0\, aq => ir23, a0 => iob23, a1 => i23, b1 => i22, b0 => iob22, bq => ir22, clk => clk3b, cq => ir21, c0 => iob21, c1 => i21, d1 => i20, d0 => iob20, dq => ir20);
  ireg_3c19 : am25s09 port map(sel => \-destimod0\, aq => ir19, a0 => iob19, a1 => i19, b1 => i18, b0 => iob18, bq => ir18, clk => clk3b, cq => ir17, c0 => iob17, c1 => i17, d1 => i16, d0 => iob16, dq => ir16);
  ireg_3d06 : am25s09 port map(sel => \-destimod1\, aq => nc371, a0 => nc372, a1 => nc373, b1 => i48, b0 => gnd, bq => ir48, clk => clk3a, cq => ir47, c0 => iob47, c1 => i47, d1 => i46, d0 => iob46, dq => ir46);
  ireg_3d07 : am25s09 port map(sel => \-destimod1\, aq => ir45, a0 => iob45, a1 => i45, b1 => i44, b0 => iob44, bq => ir44, clk => clk3a, cq => ir43, c0 => iob43, c1 => i43, d1 => i42, d0 => iob42, dq => ir42);
  ireg_3d16 : am25s09 port map(sel => \-destimod1\, aq => ir41, a0 => iob41, a1 => i41, b1 => i40, b0 => iob40, bq => ir40, clk => clk3b, cq => ir39, c0 => iob39, c1 => i39, d1 => i38, d0 => iob38, dq => ir38);
  ireg_3d17 : am25s09 port map(sel => \-destimod1\, aq => ir37, a0 => iob37, a1 => i37, b1 => i36, b0 => iob36, bq => ir36, clk => clk3b, cq => ir35, c0 => iob35, c1 => i35, d1 => i34, d0 => iob34, dq => ir34);
  ireg_3d18 : am25s09 port map(sel => \-destimod1\, aq => ir33, a0 => iob33, a1 => i33, b1 => i32, b0 => iob32, bq => ir32, clk => clk3b, cq => ir31, c0 => iob31, c1 => i31, d1 => i30, d0 => iob30, dq => ir30);
  ireg_3d19 : am25s09 port map(sel => \-destimod1\, aq => ir29, a0 => iob29, a1 => i29, b1 => i28, b0 => iob28, bq => ir28, clk => clk3b, cq => ir27, c0 => iob27, c1 => i27, d1 => i26, d0 => iob26, dq => ir26);
  ireg_3d20 : am25s09 port map(sel => \-destimod0\, aq => nc374, a0 => nc375, a1 => nc376, b1 => nc377, b0 => nc378, bq => nc379, clk => clk3b, cq => ir25, c0 => iob25, c1 => i25, d1 => i24, d0 => iob24, dq => ir24);
end architecture;
