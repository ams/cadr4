library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sip220_330_8 is
  port (
    r2 : out std_logic;
    r3 : out std_logic;
    r4 : out std_logic;
    r5 : out std_logic;
    r6 : out std_logic;
    r7 : out std_logic
    );
end;

architecture ttl of sip220_330_8 is
begin

end;
