library ieee;
use ieee.std_logic_1164.all;

entity cadr4_tb is
end;

architecture testbench of cadr4_tb is

  component cadr4 is
  end component;

begin

end;
