library ieee;
use ieee.std_logic_1164.all;

entity busint_xa is
  port (
    \-lm power reset\ : in     std_logic;
    \-xaddrdrive\   : in     std_logic;
    \xaddr par out\ : in     std_logic;
    \xbus extgrant out\ : in     std_logic;
    \xbus request\  : in     std_logic;
    clk0            : in     std_logic;
    reset           : in     std_logic;
    xao0            : in     std_logic;
    xao1            : in     std_logic;
    xao10           : in     std_logic;
    xao11           : in     std_logic;
    xao12           : in     std_logic;
    xao13           : in     std_logic;
    xao14           : in     std_logic;
    xao15           : in     std_logic;
    xao16           : in     std_logic;
    xao17           : in     std_logic;
    xao18           : in     std_logic;
    xao19           : in     std_logic;
    xao2            : in     std_logic;
    xao20           : in     std_logic;
    xao21           : in     std_logic;
    xao3            : in     std_logic;
    xao4            : in     std_logic;
    xao5            : in     std_logic;
    xao6            : in     std_logic;
    xao7            : in     std_logic;
    xao8            : in     std_logic;
    xao9            : in     std_logic;
    \-xaddr par\    : inout  std_logic;
    \-xaddr0\       : inout  std_logic;
    \-xaddr10\      : inout  std_logic;
    \-xaddr11\      : inout  std_logic;
    \-xaddr12\      : inout  std_logic;
    \-xaddr13\      : inout  std_logic;
    \-xaddr14\      : inout  std_logic;
    \-xaddr15\      : inout  std_logic;
    \-xaddr16\      : inout  std_logic;
    \-xaddr17\      : inout  std_logic;
    \-xaddr18\      : inout  std_logic;
    \-xaddr19\      : inout  std_logic;
    \-xaddr1\       : inout  std_logic;
    \-xaddr20\      : inout  std_logic;
    \-xaddr21\      : inout  std_logic;
    \-xaddr2\       : inout  std_logic;
    \-xaddr3\       : inout  std_logic;
    \-xaddr4\       : inout  std_logic;
    \-xaddr5\       : inout  std_logic;
    \-xaddr6\       : inout  std_logic;
    \-xaddr7\       : inout  std_logic;
    \-xaddr8\       : inout  std_logic;
    \-xaddr9\       : inout  std_logic;
    \-xbus ack\     : inout  std_logic;
    \-xbus busy\    : inout  std_logic;
    \-xbus extgrant out\ : inout  std_logic;
    \-xbus extrq\   : inout  std_logic;
    \-xbus init\    : inout  std_logic;
    \-xbus intr\    : inout  std_logic;
    \-xbus power reset\ : inout  std_logic;
    \-xbus rq\      : inout  std_logic;
    \-xbus sync\    : inout  std_logic;
    \lm power reset\ : out    std_logic;
    \xbus ack in\   : out    std_logic;
    \xbus busy in\  : out    std_logic;
    \xbus extrq in\ : out    std_logic;
    \xbus intr in\  : out    std_logic
  );
end entity;
