library ieee;
use ieee.std_logic_1164.all;

package unsorted is

component ic_16dummy port(dummy:in std_logic);end component;
component ic_2147 port(a0:in std_logic;a1:in std_logic;a2:in std_logic;a3:in std_logic;a4:in std_logic;a5:in std_logic;do:out std_logic;we_n:in std_logic;ce_n:in std_logic;di:in std_logic;a11:in std_logic;a10:in std_logic;a9:in std_logic;a8:in std_logic;a7:in std_logic;a6:in std_logic);end component;
component ic_2507 port(i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;i4:in std_logic;i5:in std_logic;d0:out std_logic;d1:out std_logic;d2:out std_logic;d3:out std_logic;d4:out std_logic;d5:out std_logic;clk:in std_logic;enb_n:in std_logic);end component;
component ic_2509 port(a0:in std_logic;a1:in std_logic;aq:out std_logic;b0:in std_logic;b1:in std_logic;bq:out std_logic;c0:in std_logic;c1:in std_logic;cq:out std_logic;d0:in std_logic;d1:in std_logic;dq:out std_logic;sel:in std_logic;clk:in std_logic);end component;
component ic_2510 port(i3:in std_logic;i2:in std_logic;i1:in std_logic;i0:in std_logic;i_1:in std_logic;i_2:in std_logic;i_3:in std_logic;sel1:in std_logic;sel0:in std_logic;ce_n:in std_logic;o3:out std_logic;o2:out std_logic;o1:out std_logic;o0:out std_logic);end component;
component ic_252519 port(o_enb_n:in std_logic;inv:in std_logic;i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;out_enb_n:in std_logic;clk:in std_logic;clk_enb_n:in std_logic;asyn_clr_n:in std_logic;q0a:out std_logic;q1a:out std_logic;q2a:out std_logic;q3a:out std_logic;q0b:out std_logic;q1b:out std_logic;q2b:out std_logic;q3b:out std_logic);end component;
component ic_5600 port(o7:out std_logic;o6:out std_logic;o5:out std_logic;o4:out std_logic;o3:out std_logic;o2:out std_logic;o1:out std_logic;o0:out std_logic;a4:in std_logic;a3:in std_logic;a2:in std_logic;a1:in std_logic;a0:in std_logic;ce_n:in std_logic);end component;
component ic_5610 port(o7:out std_logic;o6:out std_logic;o5:out std_logic;o4:out std_logic;o3:out std_logic;o2:out std_logic;o1:out std_logic;o0:out std_logic;a4:in std_logic;a3:in std_logic;a2:in std_logic;a1:in std_logic;a0:in std_logic;ce_n:in std_logic);end component;
component ic_7400 port(g1b:in std_logic;g1a:in std_logic;g1q_n:out std_logic;g2b:in std_logic;g2a:in std_logic;g2q_n:out std_logic;g3b:in std_logic;g3a:in std_logic;g3q_n:out std_logic;g4q_n:out std_logic;g4a:in std_logic;g4b:in std_logic);end component;
component ic_7402 port(g1q_n:out std_logic;g1a:in std_logic;g1b:in std_logic;g2q_n:out std_logic;g2a:in std_logic;g2b:in std_logic;g3b:in std_logic;g3a:in std_logic;g3q_n:out std_logic;g4b:in std_logic;g4a:in std_logic;g4q_n:out std_logic);end component;
component ic_7404 port(g1a:in std_logic;g1q_n:out std_logic;g2a:in std_logic;g2q_n:out std_logic;g3a:in std_logic;g3q_n:out std_logic;g4q:out std_logic;g4a:in std_logic;g5q_n:out std_logic;g5a:in std_logic;g6q_n:out std_logic;g6a:in std_logic);end component;
component ic_7408 port(g1b:in std_logic;g1a:in std_logic;g1q:out std_logic;g2b:in std_logic;g2a:in std_logic;g2q:out std_logic;g3a:in std_logic;g3b:in std_logic;g3q:out std_logic;g4q:out std_logic;g4a:in std_logic;g4b:in std_logic);end component;
component ic_7410 port(g1a:in std_logic;g1b:in std_logic;g2a:in std_logic;g2b:in std_logic;g2c:in std_logic;g2y_n:out std_logic;g3y_n:out std_logic;g3a:in std_logic;g3b:in std_logic;g3c:in std_logic;g1y_n:out std_logic;g1c:in std_logic);end component;
component ic_74109 port(clr1_n:in std_logic;j1:in std_logic;k1_n:in std_logic;clk1:in std_logic;pre1_n:in std_logic;q1:out std_logic;q1_n:out std_logic;clr2_n:in std_logic;j2:in std_logic;k2_n:in std_logic;clk2:in std_logic;pre2_n:in std_logic;q2:out std_logic;q2_n:out std_logic);end component;
component ic_7411 port(g1a:in std_logic;g1b:in std_logic;g2a:in std_logic;g2b:in std_logic;g2c:in std_logic;g2y_n:out std_logic;g3y_n:out std_logic;g3a:in std_logic;g3b:in std_logic;g3c:in std_logic;g1y_n:out std_logic;g1c:in std_logic);end component;
component ic_74133 port(g:in std_logic;f:in std_logic;e:in std_logic;d:in std_logic;c:in std_logic;b:in std_logic;a:in std_logic;q_n:out std_logic;h:in std_logic;i:in std_logic;j:in std_logic;k:in std_logic;l:in std_logic;m:in std_logic);end component;
component ic_74138 port(a:in std_logic;b:in std_logic;c:in std_logic;g2a:in std_logic;g2b:in std_logic;g1:in std_logic;y7:out std_logic;y6:out std_logic;y5:out std_logic;y4:out std_logic;y3:out std_logic;y2:out std_logic;y1:out std_logic;y0:out std_logic);end component;
component ic_74139 port(g1:in std_logic;a1:in std_logic;b1:in std_logic;g1y0:out std_logic;g1y1:out std_logic;g1y2:out std_logic;g1y3:out std_logic;g2y3:out std_logic;g2y2:out std_logic;g2y1:out std_logic;g2y0:out std_logic;b2:in std_logic;a2:in std_logic;g2:in std_logic);end component;
component ic_7414 port(g1a:in std_logic;g1q_n:out std_logic;g2a:in std_logic;g2q_n:out std_logic;g3a:in std_logic;g3q_n:out std_logic;g4q:out std_logic;g4a:in std_logic;g5q_n:out std_logic;g5a:in std_logic;g6q_n:out std_logic;g6a:in std_logic);end component;
component ic_74151 port(i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;i4:in std_logic;i5:in std_logic;i6:in std_logic;i7:in std_logic;q:out std_logic;q_n:out std_logic;sel2:in std_logic;sel1:in std_logic;sel0:in std_logic;ce_n:in std_logic);end component;
component ic_74153 port(enb1_n:in std_logic;sel1:in std_logic;g1c3:in std_logic;g1c2:in std_logic;g1c1:in std_logic;g1c0:in std_logic;g1q:out std_logic;g2q:out std_logic;g2c0:in std_logic;g2c1:in std_logic;g2c2:in std_logic;g2c3:in std_logic;sel0:in std_logic;enb2_n:in std_logic);end component;
component ic_74157 port(sel:in std_logic;a4:in std_logic;b4:in std_logic;y4:out std_logic;a3:in std_logic;b3:in std_logic;y3:out std_logic;y2:out std_logic;b2:in std_logic;a2:in std_logic;y1:out std_logic;b1:in std_logic;a1:in std_logic;enb_n:in std_logic);end component;
component ic_74169 port(co_n:out std_logic;i3:in std_logic;i2:in std_logic;i1:in std_logic;i0:in std_logic;o3:out std_logic;o2:out std_logic;o1:out std_logic;o0:out std_logic;enb_t_n:in std_logic;enb_p_n:in std_logic;load_n:in std_logic;up_dn:in std_logic;clk:in std_logic);end component;
component ic_74174 port(clr_n:in std_logic;q1:in std_logic;d1:in std_logic;d2:in std_logic;q2:in std_logic;d3:in std_logic;q3:in std_logic;clk:in std_logic;q4:in std_logic;d4:in std_logic;q5:in std_logic;d5:in std_logic;d6:in std_logic;q6:in std_logic);end component;
component ic_74175 port(d0:in std_logic;q0:out std_logic;q0_n:out std_logic;d1:in std_logic;q1:out std_logic;q1_n:out std_logic;d2:in std_logic;q2:out std_logic;q2_n:out std_logic;d3:in std_logic;q3:out std_logic;q3_n:out std_logic;clr_n:in std_logic;clk:in std_logic);end component;
component ic_74181 port(cout_n:out std_logic;y:out std_logic;x:out std_logic;aeb:out std_logic;f3:out std_logic;f2:out std_logic;f1:out std_logic;f0:out std_logic;b3:in std_logic;b2:in std_logic;b1:in std_logic;b0:in std_logic;a3:in std_logic;a2:in std_logic;a1:in std_logic;a0:in std_logic;m:in std_logic;s3:in std_logic;s2:in std_logic;s1:in std_logic;s0:in std_logic;cin_n:in std_logic);end component;
component ic_74182 port(xout:out std_logic;yout:out std_logic;x3:out std_logic;y3:out std_logic;cout2_n:out std_logic;x2:in std_logic;y2:in std_logic;cout1_n:out std_logic;x1:in std_logic;y1:in std_logic;cout0_n:out std_logic;x0:in std_logic;y0:in std_logic;cin_n:in std_logic);end component;
component ic_74194 port(clr_n:in std_logic;sir:in std_logic;i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;sil:in std_logic;s0:in std_logic;s1:in std_logic;clk:in std_logic;q3:out std_logic;q2:out std_logic;q1:out std_logic;q0:out std_logic);end component;
component ic_7420 port(g1a:in std_logic;g1b:in std_logic;g1c:in std_logic;g1d:in std_logic;g1y_n:out std_logic;g2y_n:out std_logic;g2a:in std_logic;g2b:in std_logic;g2c:in std_logic;g2d:in std_logic);end component;
component ic_74240 port(aenb_n:in std_logic;ain0:in std_logic;bout3:out std_logic;ain1:in std_logic;bout2:out std_logic;ain2:in std_logic;bout1:out std_logic;ain3:in std_logic;bout0:out std_logic;bin0:in std_logic;aout3:out std_logic;bin1:in std_logic;aout2:out std_logic;bin2:in std_logic;aout1:out std_logic;bin3:in std_logic;aout0:out std_logic;benb_n:in std_logic);end component;
component ic_74241 port(aenb_n:in std_logic;ain0:in std_logic;bout3:out std_logic;ain1:in std_logic;bout2:out std_logic;ain2:in std_logic;bout1:out std_logic;ain3:in std_logic;bout0:out std_logic;bin0:in std_logic;aout3:out std_logic;bin1:in std_logic;aout2:out std_logic;bin2:in std_logic;aout1:out std_logic;bin3:in std_logic;aout0:out std_logic;benb:in std_logic);end component;
component ic_74244 port(aenb_n:in std_logic;ain0:in std_logic;bout3:out std_logic;ain1:in std_logic;bout2:out std_logic;ain2:in std_logic;bout1:out std_logic;ain3:in std_logic;bout0:out std_logic;bin0:in std_logic;aout3:out std_logic;bin1:in std_logic;aout2:out std_logic;bin2:in std_logic;aout1:out std_logic;bin3:in std_logic;aout0:out std_logic;benb_n:in std_logic);end component;
component ic_74258 port(a0:in std_logic;a1:in std_logic;ay:out std_logic;b0:in std_logic;b1:in std_logic;by:out std_logic;c0:in std_logic;c1:in std_logic;cy:out std_logic;d0:in std_logic;d1:in std_logic;dy:out std_logic;sel:in std_logic;enb_n:in std_logic);end component;
component ic_74260 port(i1:in std_logic;i2:in std_logic;i3:in std_logic;o1:out std_logic;i4:in std_logic;i5:in std_logic);end component;
component ic_7428 port(g1q_n:out std_logic;g1a:in std_logic;g1b:in std_logic;g2q_n:out std_logic;g2a:in std_logic;g2b:in std_logic;g3a:in std_logic;g3b:in std_logic;g3q_n:out std_logic;g4a:in std_logic;g4b:in std_logic;g4q_n:out std_logic);end component;
component ic_74280 port(i0:in std_logic;i1:in std_logic;i2:in std_logic;even:out std_logic;odd:out std_logic;i3:in std_logic;i4:in std_logic;i5:in std_logic;i6:in std_logic;i7:in std_logic;i8:in std_logic);end component;
component ic_74283 port(c4:out std_logic;a3:in std_logic;a2:in std_logic;a1:in std_logic;a0:in std_logic;s3:out std_logic;s2:out std_logic;s1:out std_logic;s0:out std_logic;b3:in std_logic;b2:in std_logic;b1:in std_logic;b0:in std_logic;c0:in std_logic);end component;
component ic_7432 port(g1a:in std_logic;g1b:in std_logic;g1y:out std_logic;g2a:in std_logic;g2b:in std_logic;g2y:out std_logic;g3y:out std_logic;g3a:in std_logic;g3b:in std_logic;g4y:out std_logic;g4a:in std_logic;g4b:in std_logic);end component;
component ic_7437 port(g1a:in std_logic;g1b:in std_logic;g1y:out std_logic;g2a:in std_logic;g2b:in std_logic;g2y:out std_logic;g3y:out std_logic;g3a:in std_logic;g3b:in std_logic;g4y:out std_logic;g4a:in std_logic;g4b:in std_logic);end component;
component ic_74373 port(i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;i4:in std_logic;i5:in std_logic;i6:in std_logic;i7:in std_logic;o0:out std_logic;o1:out std_logic;o2:out std_logic;o3:out std_logic;o4:out std_logic;o5:out std_logic;o6:out std_logic;o7:out std_logic;hold_n:in std_logic;oenb_n:in std_logic);end component;
component ic_74374 port(i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;i4:in std_logic;i5:in std_logic;i6:in std_logic;i7:in std_logic;o0:out std_logic;o1:out std_logic;o2:out std_logic;o3:out std_logic;o4:out std_logic;o5:out std_logic;o6:out std_logic;o7:out std_logic;clk:in std_logic;oenb_n:in std_logic);end component;
component ic_74472 port(a0:in std_logic;a1:in std_logic;a2:in std_logic;a3:in std_logic;a4:in std_logic;d0:in std_logic;d1:in std_logic;d2:in std_logic;d3:in std_logic;d4:in std_logic;d5:in std_logic;d6:in std_logic;d7:in std_logic;ce_n:in std_logic;a5:in std_logic;a6:in std_logic;a7:in std_logic;a8:in std_logic);end component;
component ic_7451 port(g1a:in std_logic;g2a:in std_logic;g2b:in std_logic;g2c:in std_logic;g2d:in std_logic;g2y:out std_logic;g1y:out std_logic;g1c:in std_logic;g1d:in std_logic;g1b:in std_logic);end component;
component ic_7464 port(d4:in std_logic;b2:in std_logic;a2:in std_logic;c3:in std_logic;b3:in std_logic;a3:in std_logic;\out\:out std_logic;a1:in std_logic;b1:in std_logic;c4:in std_logic;b4:in std_logic;a4:in std_logic);end component;
component ic_7474 port(g1r_n:in std_logic;g1d:in std_logic;g1clk:in std_logic;g1s_n:in std_logic;g1q:out std_logic;g1q_n:out std_logic;g2q_n:out std_logic;g2q:out std_logic;g2s_n:in std_logic;g2clk:in std_logic;g2d:in std_logic;g2r_n:in std_logic);end component;
component ic_7486 port(g1a:in std_logic;g1b:in std_logic;g1y:out std_logic;g2a:in std_logic;g2b:in std_logic;g2y:out std_logic;g3y:out std_logic;g3a:in std_logic;g3b:in std_logic;g4y:out std_logic;g4a:in std_logic;g4b:in std_logic);end component;
component ic_8221 port(d1:out std_logic;i1:in std_logic;we1_n:in std_logic;i0:in std_logic;d0:out std_logic;we0_n:in std_logic;a0:in std_logic;a1:in std_logic;a2:in std_logic;a3:in std_logic;a4:in std_logic;strobe:in std_logic;wclk_n:in std_logic;ce:in std_logic);end component;
component ic_9328 port(clr_n:in std_logic;aq_n:in std_logic;aq:in std_logic;asel:in std_logic;ai1:in std_logic;ai0:in std_logic;aclk:in std_logic;comclk:in std_logic;bclk:in std_logic;bi0:in std_logic;bi1:in std_logic;bsel:in std_logic;bq:in std_logic;bq_n:in std_logic);end component;
component ic_93425a port(a0:in std_logic;a1:in std_logic;a2:in std_logic;a3:in std_logic;a4:in std_logic;a5:in std_logic;a6:in std_logic;a7:in std_logic;a8:in std_logic;a9:in std_logic;ce_n:in std_logic;we_n:in std_logic;di:in std_logic;do:out std_logic);end component;
component ic_9346 port(a5:in std_logic;a4:in std_logic;a3:in std_logic;a2:in std_logic;a1:in std_logic;a0:in std_logic;b5:in std_logic;b4:in std_logic;b3:in std_logic;b2:in std_logic;b1:in std_logic;b0:in std_logic;enb:in std_logic;eq:out std_logic);end component;
component ic_9348 port(i0:in std_logic;i1:in std_logic;i2:in std_logic;i3:in std_logic;i4:in std_logic;i5:in std_logic;i6:in std_logic;i7:in std_logic;i8:in std_logic;i9:in std_logic;i10:in std_logic;i11:in std_logic;pe:out std_logic;po:out std_logic);end component;
component ic_942_1 port(g1a1:in std_logic;g1b1:in std_logic;g2a1:in std_logic;g2b1:in std_logic;g2c1:in std_logic;g2d1:in std_logic;out1:out std_logic;g1a2:in std_logic;g1b2:in std_logic;g2a2:in std_logic;g2b2:in std_logic;g2c2:in std_logic;g2d2:in std_logic;out2:out std_logic);end component;
component ic_res20 port(r2:in std_logic;r3:in std_logic;r4:in std_logic;r5:in std_logic;r6:in std_logic;r7:in std_logic;r8:in std_logic;r9:in std_logic;r10:in std_logic;r11:in std_logic;r12:in std_logic;r13:in std_logic;r14:in std_logic;r15:in std_logic;r16:in std_logic;r17:in std_logic;r18:in std_logic;r19:in std_logic);end component;
component ic_sip220_330_8 port(r2:in std_logic;r3:in std_logic;r4:in std_logic;r5:in std_logic;r6:in std_logic;r7:in std_logic);end component;
component ic_sip330_470_8 port(r2:in std_logic;r3:in std_logic;r4:in std_logic;r5:in std_logic;r6:in std_logic;r7:in std_logic);end component;
component ic_td100 port(input:in std_logic;o_20ns:out std_logic;o_40ns:out std_logic;o_60ns:out std_logic;o_80ns:out std_logic;o_100ns:out std_logic);end component;
component ic_td25 port(input:in std_logic;o_10ns:out std_logic;o_20ns:out std_logic;o_25ns:out std_logic;o_15ns:out std_logic;o_5ns:out std_logic);end component;
component ic_td250 port(input:in std_logic;o_50ns:out std_logic;o_100ns:out std_logic;o_150ns:out std_logic;o_200ns:out std_logic;o_250ns:out std_logic);end component;
component ic_td50 port(input:in std_logic;o_10ns:out std_logic;o_20ns:out std_logic;o_30ns:out std_logic;o_40ns:out std_logic;o_50ns:out std_logic);end component;
component ic_til309 port(l2:in std_logic;l4:in std_logic;l8:in std_logic;l1:in std_logic;latch:in std_logic;i4:in std_logic;i8:in std_logic;i2:in std_logic;blank_n:in std_logic;dp:in std_logic;test_n:in std_logic;ldp:in std_logic;i1:in std_logic);end component;

alias ic_25ls2519 is ic_252519;
alias ic_25s07 is ic_2507;
alias ic_25s09 is ic_2509;
alias ic_25s10 is ic_2510;
alias ic_74ls109 is ic_74109;
alias ic_74ls14 is ic_7414;
alias ic_74ls244 is ic_74244;
alias ic_74s00 is ic_7400;
alias ic_74s02 is ic_7402;
alias ic_74s04 is ic_7404;
alias ic_74s08 is ic_7408;
alias ic_74s10 is ic_7410;
alias ic_74s11 is ic_7411;
alias ic_74s133 is ic_74133;
alias ic_74s138 is ic_74138;
alias ic_74s139 is ic_74139;
alias ic_74s151 is ic_74151;
alias ic_74s153 is ic_74153;
alias ic_74s157 is ic_74157;
alias ic_74s169 is ic_74169;
alias ic_74s174 is ic_74174;
alias ic_74s175 is ic_74175;
alias ic_74s181 is ic_74181;
alias ic_74s182 is ic_74182;
alias ic_74s194 is ic_74194;
alias ic_74s20 is ic_7420;
alias ic_74s240 is ic_74240;
alias ic_74s241 is ic_74241;
alias ic_74s258 is ic_74258;
alias ic_74s260 is ic_74260;
alias ic_74s280 is ic_74280;
alias ic_74s283 is ic_74283;
alias ic_74s32 is ic_7432;
alias ic_74s37 is ic_7437;
alias ic_74s373 is ic_74373;
alias ic_74s374 is ic_74374;
alias ic_74s472 is ic_74472;
alias ic_74s51 is ic_7451;
alias ic_74s64 is ic_7464;
alias ic_74s74 is ic_7474;
alias ic_74s86 is ic_7486;
alias ic_82s21 is ic_8221;
alias ic_93s46 is ic_9346;
alias ic_93s48 is ic_9348;
alias ic_9s42_1 is ic_942_1;

end;

package body unsorted is

end;
