library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_pdlctl is
  port (
    \-reset\      : in  std_logic;
    pdlwrited     : out std_logic;
    \-pdlwrited\  : out std_logic;
    pdlwrite      : out std_logic;
    \-destpdl(x)\ : in  std_logic;
    pwidx         : out std_logic;
    \-pwidx\      : out std_logic;
    clk4f         : in  std_logic;
    imodd         : out std_logic;
    \-imodd\      : out std_logic;
    imod          : in  std_logic;
    \-destspc\    : in  std_logic;
    \-destspcd\   : out std_logic;
    \-pdlpb\      : out std_logic;
    pdlptr0       : in  std_logic;
    pdlidx0       : in  std_logic;
    \-pdla0b\     : out std_logic;
    pdlptr1       : in  std_logic;
    pdlidx1       : in  std_logic;
    \-pdla1b\     : out std_logic;
    \-pdla2b\     : out std_logic;
    pdlidx2       : in  std_logic;
    pdlptr2       : in  std_logic;
    \-pdla3b\     : out std_logic;
    pdlidx3       : in  std_logic;
    pdlptr3       : in  std_logic;
    gnd           : in  std_logic;
    \-pdlpa\      : out std_logic;
    pdlptr8       : in  std_logic;
    pdlidx8       : in  std_logic;
    \-pdla8b\     : out std_logic;
    pdlptr9       : in  std_logic;
    pdlidx9       : in  std_logic;
    \-pdla9b\     : out std_logic;
    \-pdla0a\     : out std_logic;
    \-pdla1a\     : out std_logic;
    \-pdla2a\     : out std_logic;
    \-pdla3a\     : out std_logic;
    \-pdla4a\     : out std_logic;
    pdlidx4       : in  std_logic;
    pdlptr4       : in  std_logic;
    \-pdla5a\     : out std_logic;
    pdlidx5       : in  std_logic;
    pdlptr5       : in  std_logic;
    \-destpdl(p)\ : in  std_logic;
    \-pdlcnt\     : out std_logic;
    clk4b         : in  std_logic;
    ir30          : in  std_logic;
    \-clk4e\      : in  std_logic;
    \-srcpdlpop\  : in  std_logic;
    \-srcpdltop\  : in  std_logic;
    pdlenb        : out std_logic;
    tse4b         : in  std_logic;
    \-pdldrive\   : out std_logic;
    \-destpdltop\ : in  std_logic;
    \-pdla4b\     : out std_logic;
    \-pdla5b\     : out std_logic;
    \-pdla6b\     : out std_logic;
    pdlidx6       : in  std_logic;
    pdlptr6       : in  std_logic;
    \-pdla7b\     : out std_logic;
    pdlidx7       : in  std_logic;
    pdlptr7       : in  std_logic;
    wp4a          : in  std_logic;
    \-pwpa\       : out std_logic;
    \-pwpb\       : out std_logic;
    \-pwpc\       : out std_logic;
    \-pdla6a\     : out std_logic;
    \-pdla7a\     : out std_logic;
    \-pdla8a\     : out std_logic;
    \-pdla9a\     : out std_logic;
    nop           : in  std_logic);
end;

architecture ttl of cadr4_pdlctl is
  signal internal19 : std_logic;
  signal nc242      : std_logic;
begin
  pdlctl_4c11 : sn74s175 port map(clr_n => \-reset\, q0 => pdlwrited, q0_n => \-pdlwrited\, d0 => pdlwrite, d1 => \-destpdl(x)\, q1_n => pwidx, q1 => \-pwidx\, clk => clk4f, q2 => imodd, q2_n => \-imodd\, d2 => imod, d3 => \-destspc\, q3_n => nc242, q3 => \-destspcd\);
  pdlctl_4c12 : sn74s258 port map(sel   => \-pdlpb\, d0 => pdlptr0, d1 => pdlidx0, dy => \-pdla0b\, c0 => pdlptr1, c1 => pdlidx1, cy => \-pdla1b\, by => \-pdla2b\, b1 => pdlidx2, b0 => pdlptr2, ay => \-pdla3b\, a1 => pdlidx3, a0 => pdlptr3, enb_n => gnd);
  pdlctl_4c16 : sn74s258 port map(sel   => \-pdlpa\, d0 => pdlptr8, d1 => pdlidx8, dy => \-pdla8b\, c0 => pdlptr9, c1 => pdlidx9, cy => \-pdla9b\, by => \-pdla0a\, b1 => pdlidx0, b0 => pdlptr0, ay => \-pdla1a\, a1 => pdlidx1, a0 => pdlptr1, enb_n => gnd);
  pdlctl_4c22 : sn74s258 port map(sel   => \-pdlpa\, d0 => pdlptr2, d1 => pdlidx2, dy => \-pdla2a\, c0 => pdlptr3, c1 => pdlidx3, cy => \-pdla3a\, by => \-pdla4a\, b1 => pdlidx4, b0 => pdlptr4, ay => \-pdla5a\, a1 => pdlidx5, a0 => pdlptr5, enb_n => gnd);
  pdlctl_4d06 : sn74s08 port map(g2b    => internal19, g2a => \-destpdl(p)\, g2q => \-pdlcnt\, g1b => '0', g1a => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  pdlctl_4d07 : sn74s51 port map(g1a    => \-pwidx\, g2a => clk4b, g2b => ir30, g2c => \-clk4e\, g2d => \-pwidx\, g2y => \-pdlpa\, g1y => \-pdlpb\, g1c => clk4b, g1d => ir30, g1b => \-clk4e\);
  pdlctl_4d08 : sn74s00 port map(g1b    => \-srcpdlpop\, g1a => \-srcpdltop\, g1q_n => pdlenb, g2b => pdlenb, g2a => tse4b, g2q_n => \-pdldrive\, g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  pdlctl_4d10 : sn74s10 port map(g1a    => \-destpdltop\, g1b => \-destpdl(x)\, g1y_n => pdlwrite, g1c => \-destpdl(p)\, g2a => '0', g2b => '0', g2c => '0', g3a => '0', g3b => '0', g3c => '0');
  pdlctl_4d14 : sn74s258 port map(sel   => \-pdlpb\, d0 => pdlptr4, d1 => pdlidx4, dy => \-pdla4b\, c0 => pdlptr5, c1 => pdlidx5, cy => \-pdla5b\, by => \-pdla6b\, b1 => pdlidx6, b0 => pdlptr6, ay => \-pdla7b\, a1 => pdlidx7, a0 => pdlptr7, enb_n => gnd);
  pdlctl_4d20 : sn74s37 port map(g1a    => pdlwrited, g1b => wp4a, g1y => \-pwpa\, g2a => pdlwrited, g2b => wp4a, g2y => \-pwpb\, g3y => \-pwpc\, g3a => wp4a, g3b => pdlwrited, g4a => '0', g4b => '0');
  pdlctl_4d24 : sn74s258 port map(sel   => \-pdlpa\, d0 => pdlptr6, d1 => pdlidx6, dy => \-pdla6a\, c0 => pdlptr7, c1 => pdlidx7, cy => \-pdla7a\, by => \-pdla8a\, b1 => pdlidx8, b0 => pdlptr8, ay => \-pdla9a\, a1 => pdlidx9, a0 => pdlptr9, enb_n => gnd);
  pdlctl_4e03 : sn74s32 port map(g3y    => internal19, g3a => \-srcpdlpop\, g3b => nop, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4a => '0', g4b => '0');
end architecture;
