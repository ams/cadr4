library ieee;
use ieee.std_logic_1164.all;

entity cadr_dram0 is
  port (
    \-dmapbenb\     : in     std_logic;
    aa0             : in     std_logic;
    aa1             : in     std_logic;
    aa2             : in     std_logic;
    aa3             : in     std_logic;
    aa4             : in     std_logic;
    aa5             : in     std_logic;
    dispwr          : in     std_logic;
    dmask0          : in     std_logic;
    dmask1          : in     std_logic;
    dmask2          : in     std_logic;
    dmask3          : in     std_logic;
    dmask4          : in     std_logic;
    dmask5          : in     std_logic;
    dmask6          : in     std_logic;
    hi4             : in     std_logic;
    hi6             : in     std_logic;
    ir12            : in     std_logic;
    ir13            : in     std_logic;
    ir14            : in     std_logic;
    ir15            : in     std_logic;
    ir16            : in     std_logic;
    ir17            : in     std_logic;
    ir18            : in     std_logic;
    ir19            : in     std_logic;
    ir20b           : in     std_logic;
    ir21b           : in     std_logic;
    ir22b           : in     std_logic;
    ir8b            : in     std_logic;
    ir9b            : in     std_logic;
    r0              : in     std_logic;
    r1              : in     std_logic;
    r2              : in     std_logic;
    r3              : in     std_logic;
    r4              : in     std_logic;
    r5              : in     std_logic;
    r6              : in     std_logic;
    vmo18           : in     std_logic;
    vmo19           : in     std_logic;
    wp2             : in     std_logic;
    \-dadr0a\       : out    std_logic;
    \-dadr10a\      : out    std_logic;
    \-dadr1a\       : out    std_logic;
    \-dadr2a\       : out    std_logic;
    \-dadr3a\       : out    std_logic;
    \-dadr4a\       : out    std_logic;
    \-dadr5a\       : out    std_logic;
    \-dadr6a\       : out    std_logic;
    \-dadr7a\       : out    std_logic;
    \-dadr8a\       : out    std_logic;
    \-dadr9a\       : out    std_logic;
    \-dwea\         : out    std_logic;
    dadr10a         : out    std_logic;
    dpc0            : out    std_logic;
    dpc1            : out    std_logic;
    dpc2            : out    std_logic;
    dpc3            : out    std_logic;
    dpc4            : out    std_logic;
    dpc5            : out    std_logic;
    ir12b           : out    std_logic;
    ir13b           : out    std_logic;
    ir14b           : out    std_logic;
    ir15b           : out    std_logic;
    ir16b           : out    std_logic;
    ir17b           : out    std_logic;
    ir18b           : out    std_logic;
    ir19b           : out    std_logic
  );
end entity cadr_dram0;
