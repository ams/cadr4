library ieee;
use ieee.std_logic_1164.all;

entity cadr_lpc is
  port (
    \lpc.hold\      : in     std_logic;
    clk4b           : in     std_logic;
    hi5             : in     std_logic;
    ir25            : in     std_logic;
    irdisp          : in     std_logic;
    pc0             : in     std_logic;
    pc1             : in     std_logic;
    pc10            : in     std_logic;
    pc11            : in     std_logic;
    pc12            : in     std_logic;
    pc13            : in     std_logic;
    pc2             : in     std_logic;
    pc3             : in     std_logic;
    pc4             : in     std_logic;
    pc5             : in     std_logic;
    pc6             : in     std_logic;
    pc7             : in     std_logic;
    pc8             : in     std_logic;
    pc9             : in     std_logic;
    lpc0            : out    std_logic;
    lpc1            : out    std_logic;
    lpc10           : out    std_logic;
    lpc11           : out    std_logic;
    lpc12           : out    std_logic;
    lpc13           : out    std_logic;
    lpc2            : out    std_logic;
    lpc3            : out    std_logic;
    lpc4            : out    std_logic;
    lpc5            : out    std_logic;
    lpc6            : out    std_logic;
    lpc7            : out    std_logic;
    lpc8            : out    std_logic;
    lpc9            : out    std_logic;
    pc0b            : out    std_logic;
    pc10b           : out    std_logic;
    pc11b           : out    std_logic;
    pc12b           : out    std_logic;
    pc13b           : out    std_logic;
    pc1b            : out    std_logic;
    pc2b            : out    std_logic;
    pc3b            : out    std_logic;
    pc4b            : out    std_logic;
    pc5b            : out    std_logic;
    pc6b            : out    std_logic;
    pc7b            : out    std_logic;
    pc8b            : out    std_logic;
    pc9b            : out    std_logic;
    wpc0            : out    std_logic;
    wpc1            : out    std_logic;
    wpc10           : out    std_logic;
    wpc11           : out    std_logic;
    wpc12           : out    std_logic;
    wpc13           : out    std_logic;
    wpc2            : out    std_logic;
    wpc3            : out    std_logic;
    wpc4            : out    std_logic;
    wpc5            : out    std_logic;
    wpc6            : out    std_logic;
    wpc7            : out    std_logic;
    wpc8            : out    std_logic;
    wpc9            : out    std_logic
  );
end entity;
