-- The MIT CADR

library ieee;
use ieee.std_logic_1164.all;

use std.env.finish;

library work;
use work.cadr_book.cadr_clockd;
use work.icmem_book.cadr_clock1;
use work.icmem_book.cadr_clock2;

entity clkgen_tb is
end;

architecture structural of clkgen_tb is

  -- clock 1 inputs

  signal \-clock reset b\ : std_logic;
  signal \-hang\          : std_logic;
  signal \-ilong\         : std_logic;
  signal gnd              : std_logic;
  signal sspeed0          : std_logic;
  signal sspeed1          : std_logic;

  -- clock 1 outputs

  signal \-tpr0\          : std_logic;
  signal \-tpr100\        : std_logic;
  signal \-tpr105\        : std_logic;
  signal \-tpr10\         : std_logic;
  signal \-tpr110\        : std_logic;
  signal \-tpr115\        : std_logic;
  signal \-tpr120\        : std_logic;
  signal \-tpr120a\       : std_logic;
  signal \-tpr125\        : std_logic;
  signal \-tpr140\        : std_logic;
  signal \-tpr15\         : std_logic;
  signal \-tpr160\        : std_logic;
  signal \-tpr180\        : std_logic;
  signal \-tpr200\        : std_logic;
  signal \-tpr20\         : std_logic;
  signal \-tpr20a\        : std_logic;
  signal \-tpr25\         : std_logic;
  signal \-tpr40\         : std_logic;
  signal \-tpr5\          : std_logic;
  signal \-tpr60\         : std_logic;
  signal \-tpr65\         : std_logic;
  signal \-tpr70\         : std_logic;
  signal \-tpr75\         : std_logic;
  signal \-tpr80\         : std_logic;
  signal \-tpr80a\        : std_logic;
  signal \-tpr85\         : std_logic;
  signal \-tprend\        : std_logic;
  signal \-tpw10\         : std_logic;
  signal \-tpw20\         : std_logic;
  signal \-tpw25\         : std_logic;
  signal \-tpw30\         : std_logic;
  signal \-tpw30a\        : std_logic;
  signal \-tpw35\         : std_logic;
  signal \-tpw40\         : std_logic;
  signal \-tpw40a\        : std_logic;
  signal \-tpw45\         : std_logic;
  signal \-tpw50\         : std_logic;
  signal \-tpw55\         : std_logic;
  signal \-tpw60\         : std_logic;
  signal \-tpw65\         : std_logic;
  signal \-tpw70\         : std_logic;
  signal \-tpw75\         : std_logic;
  signal cyclecompleted   : std_logic;  
  signal tprend           : std_logic;
  
  -- clock 2 inputs

  signal \machruna l\     : std_logic;
  signal machrun          : std_logic;
  signal hi1              : std_logic;

  -- clock 2 outputs

  signal clk4             : std_logic;
  signal \-clk0\          : std_logic;
  signal mclk7            : std_logic;
  signal \-mclk0\         : std_logic;
  signal \-wp1\           : std_logic;
  signal tpwp             : std_logic;
  signal \-wp2\           : std_logic;
  signal \-wp3\           : std_logic;
  signal \-wp4\           : std_logic;
  signal tpclk            : std_logic;
  signal \-tptse\         : std_logic;
  signal \-tpclk\         : std_logic;
  signal tptse            : std_logic;  
  signal tpwpiram         : std_logic;
  signal \-wp5\           : std_logic;
  signal clk5             : std_logic;
  signal mclk5            : std_logic;
  signal \-tse1\          : std_logic;
  signal \-tse2\          : std_logic;
  signal \-tse3\          : std_logic;
  signal \-tse4\          : std_logic;
  signal clk1             : std_logic;
  signal clk2             : std_logic;
  signal clk3             : std_logic;
  signal mclk1            : std_logic;
  
  -- clockd inputs
  
  signal reset          : std_logic;
  signal hi2            : std_logic;
  signal hi3            : std_logic;
  signal hi4            : std_logic;
  signal hi5            : std_logic;
  signal hi6            : std_logic;
  signal hi7            : std_logic;
  signal hi8            : std_logic;
  signal hi9            : std_logic;
  signal hi10           : std_logic;
  signal hi11           : std_logic;
  signal hi12           : std_logic;
  signal lcry3          : std_logic;
  signal \-srcpdlptr\   : std_logic;
  signal \-srcpdlidx\   : std_logic;

  -- clockd outputs

  signal \-clk1\        : std_logic;
  signal clk1a          : std_logic;
  signal \-reset\       : std_logic;
  signal mclk1a         : std_logic;
  signal \-mclk1\       : std_logic;
  signal wp1b           : std_logic;
  signal wp1a           : std_logic;
  signal tse1b          : std_logic;
  signal tse1a          : std_logic;
  signal \-upperhighok\ : std_logic;
  signal \-lcry3\       : std_logic;
  signal \-clk2c\       : std_logic;
  signal \-clk2a\       : std_logic;
  signal wp2            : std_logic;
  signal tse2           : std_logic;
  signal clk2a          : std_logic;
  signal clk2b          : std_logic;
  signal clk2c          : std_logic;
  signal \-clk3a\       : std_logic;
  signal clk3a          : std_logic;
  signal clk3b          : std_logic;
  signal clk3c          : std_logic;
  signal \-clk3g\       : std_logic;
  signal \-clk3d\       : std_logic;
  signal wp3a           : std_logic;
  signal tse3a          : std_logic;
  signal clk3d          : std_logic;
  signal clk3e          : std_logic;
  signal clk3f          : std_logic;
  signal \-clk4a\       : std_logic;
  signal clk4a          : std_logic;
  signal clk4b          : std_logic;
  signal clk4c          : std_logic;
  signal \-clk4e\       : std_logic;
  signal \-clk4d\       : std_logic;
  signal wp4c           : std_logic;
  signal wp4b           : std_logic;
  signal wp4a           : std_logic;
  signal clk4d          : std_logic;
  signal clk4e          : std_logic;
  signal clk4f          : std_logic;
  signal tse4b          : std_logic;
  signal tse4a          : std_logic;
  signal srcpdlptr      : std_logic;
  signal srcpdlidx      : std_logic;

begin

  --- Clock Generation (clkgen)
  i_clock1 : entity work.cadr_clock1(mete) port map(\-clock reset b\ => \-clock reset b\, \-hang\ => \-hang\, cyclecompleted => cyclecompleted, \-tpr0\ => \-tpr0\, \-tpr40\ => \-tpr40\, gnd => gnd, \-tprend\ => \-tprend\, \-tpw20\ => \-tpw20\, \-tpw40\ => \-tpw40\, \-tpw50\ => \-tpw50\, \-tpw30\ => \-tpw30\, \-tpw10\ => \-tpw10\, \-tpw60\ => \-tpw60\, \-tpw70\ => \-tpw70\, \-tpw75\ => \-tpw75\, \-tpw65\ => \-tpw65\, \-tpw55\ => \-tpw55\, \-tpw30a\ => \-tpw30a\, \-tpw40a\ => \-tpw40a\, \-tpw45\ => \-tpw45\, \-tpw35\ => \-tpw35\, \-tpw25\ => \-tpw25\, \-tpr100\ => \-tpr100\, \-tpr140\ => \-tpr140\, \-tpr160\ => \-tpr160\, tprend => tprend, sspeed1 => sspeed1, sspeed0 => sspeed0, \-ilong\ => \-ilong\, \-tpr75\ => \-tpr75\, \-tpr115\ => \-tpr115\, \-tpr85\ => \-tpr85\, \-tpr125\ => \-tpr125\, \-tpr10\ => \-tpr10\, \-tpr20a\ => \-tpr20a\, \-tpr25\ => \-tpr25\, \-tpr15\ => \-tpr15\, \-tpr5\ => \-tpr5\, \-tpr80\ => \-tpr80\, \-tpr60\ => \-tpr60\, \-tpr20\ => \-tpr20\, \-tpr180\ => \-tpr180\, \-tpr200\ => \-tpr200\, \-tpr120\ => \-tpr120\, \-tpr110\ => \-tpr110\, \-tpr120a\ => \-tpr120a\, \-tpr105\ => \-tpr105\, \-tpr70\ => \-tpr70\, \-tpr80a\ => \-tpr80a\, \-tpr65\ => \-tpr65\);
  i_clock2 : entity work.cadr_clock2(mete) port map(clk4 => clk4, \-clk0\ => \-clk0\, gnd => gnd, mclk7 => mclk7, \-mclk0\ => \-mclk0\, \-wp1\ => \-wp1\, tpwp => tpwp, \-wp2\ => \-wp2\, \-wp3\ => \-wp3\, \-wp4\ => \-wp4\, \-tprend\ => \-tprend\, tpclk => tpclk, \-tptse\ => \-tptse\, \-tpr25\ => \-tpr25\, \-clock reset b\ => \-clock reset b\, tptse => tptse, \-tpw70\ => \-tpw70\, \-tpclk\ => \-tpclk\, \-tpr0\ => \-tpr0\, \-tpr5\ => \-tpr5\, \-tpw30\ => \-tpw30\, \machruna l\ => \machruna l\, tpwpiram => tpwpiram, \-wp5\ => \-wp5\, clk5 => clk5, mclk5 => mclk5, \-tpw45\ => \-tpw45\, \-tse1\ => \-tse1\, \-tse2\ => \-tse2\, \-tse3\ => \-tse3\, \-tse4\ => \-tse4\, clk1 => clk1, clk2 => clk2, clk3 => clk3, mclk1 => mclk1, machrun => machrun, hi1 => hi1);
  i_clockd : cadr_clockd port map(\-clk1\ => \-clk1\, hi12 => hi12, clk1a => clk1a, reset => reset, \-reset\ => \-reset\, mclk1a => mclk1a, \-mclk1\ => \-mclk1\, mclk1 => mclk1, clk1 => clk1, \-wp1\ => \-wp1\, wp1b => wp1b, wp1a => wp1a, tse1b => tse1b, \-tse1\ => \-tse1\, tse1a => tse1a, hi1 => hi1, hi2 => hi2, hi3 => hi3, hi4 => hi4, hi5 => hi5, hi6 => hi6, hi7 => hi7, \-upperhighok\ => \-upperhighok\, hi8 => hi8, hi9 => hi9, hi10 => hi10, hi11 => hi11, lcry3 => lcry3, \-lcry3\ => \-lcry3\, clk2 => clk2, \-clk2c\ => \-clk2c\, \-clk2a\ => \-clk2a\, wp2 => wp2, \-wp2\ => \-wp2\, tse2 => tse2, \-tse2\ => \-tse2\, clk2a => clk2a, clk2b => clk2b, clk2c => clk2c, \-clk3a\ => \-clk3a\, clk3a => clk3a, clk3b => clk3b, clk3c => clk3c, clk3 => clk3, \-clk3g\ => \-clk3g\, \-clk3d\ => \-clk3d\, wp3a => wp3a, \-wp3\ => \-wp3\, tse3a => tse3a, \-tse3\ => \-tse3\, clk3d => clk3d, clk3e => clk3e, clk3f => clk3f, \-clk4a\ => \-clk4a\, clk4a => clk4a, clk4b => clk4b, clk4c => clk4c, clk4 => clk4, \-clk4e\ => \-clk4e\, \-clk4d\ => \-clk4d\, wp4c => wp4c, \-wp4\ => \-wp4\, wp4b => wp4b, wp4a => wp4a, clk4d => clk4d, clk4e => clk4e, clk4f => clk4f, \-tse4\ => \-tse4\, tse4b => tse4b, tse4a => tse4a, srcpdlptr => srcpdlptr, \-srcpdlptr\ => \-srcpdlptr\, srcpdlidx => srcpdlidx, \-srcpdlidx\ => \-srcpdlidx\);

  -- fixed inputs, minimum speed=00, no long instruction, no hang

  -- clock1
  gnd       <= '0';
  sspeed1   <= '0';
  sspeed0   <= '1';
  \-ilong\  <= not '0';
  \-hang\   <= not '0';

  -- clock2
  hi1          <= '1';
  machrun      <= '1';
  \machruna l\ <= not machrun; -- -machrun

  -- clockd
  reset          <= not \-clock reset b\;
  hi2            <= '1';
  hi3            <= '1';
  hi4            <= '1';
  hi5            <= '1';
  hi6            <= '1';
  hi7            <= '1';
  hi8            <= '1';
  hi9            <= '1';
  hi10           <= '1';
  hi11           <= '1';
  hi12           <= '1';
  lcry3          <= '0';
  \-srcpdlptr\   <= '0';
  \-srcpdlidx\   <= '0';

  process
  begin
    \-clock reset b\ <= '0';
    wait for 10 ns;
    \-clock reset b\ <= not '0';
    wait for 1000 ns;
    finish;
  end process;

end architecture;
