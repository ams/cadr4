library ieee;
use ieee.std_logic_1164.all;

entity cadr_ireg is
  port (
    \-destimod0\    : in     std_logic;
    \-destimod1\    : in     std_logic;
    clk3a           : in     std_logic;
    clk3b           : in     std_logic;
    i0              : in     std_logic;
    i1              : in     std_logic;
    i10             : in     std_logic;
    i11             : in     std_logic;
    i12             : in     std_logic;
    i13             : in     std_logic;
    i14             : in     std_logic;
    i15             : in     std_logic;
    i16             : in     std_logic;
    i17             : in     std_logic;
    i18             : in     std_logic;
    i19             : in     std_logic;
    i2              : in     std_logic;
    i20             : in     std_logic;
    i21             : in     std_logic;
    i22             : in     std_logic;
    i23             : in     std_logic;
    i24             : in     std_logic;
    i25             : in     std_logic;
    i26             : in     std_logic;
    i27             : in     std_logic;
    i28             : in     std_logic;
    i29             : in     std_logic;
    i3              : in     std_logic;
    i30             : in     std_logic;
    i31             : in     std_logic;
    i32             : in     std_logic;
    i33             : in     std_logic;
    i34             : in     std_logic;
    i35             : in     std_logic;
    i36             : in     std_logic;
    i37             : in     std_logic;
    i38             : in     std_logic;
    i39             : in     std_logic;
    i4              : in     std_logic;
    i40             : in     std_logic;
    i41             : in     std_logic;
    i42             : in     std_logic;
    i43             : in     std_logic;
    i44             : in     std_logic;
    i45             : in     std_logic;
    i46             : in     std_logic;
    i47             : in     std_logic;
    i48             : in     std_logic;
    i5              : in     std_logic;
    i6              : in     std_logic;
    i7              : in     std_logic;
    i8              : in     std_logic;
    i9              : in     std_logic;
    iob0            : in     std_logic;
    iob1            : in     std_logic;
    iob10           : in     std_logic;
    iob11           : in     std_logic;
    iob12           : in     std_logic;
    iob13           : in     std_logic;
    iob14           : in     std_logic;
    iob15           : in     std_logic;
    iob16           : in     std_logic;
    iob17           : in     std_logic;
    iob18           : in     std_logic;
    iob19           : in     std_logic;
    iob2            : in     std_logic;
    iob20           : in     std_logic;
    iob21           : in     std_logic;
    iob22           : in     std_logic;
    iob23           : in     std_logic;
    iob24           : in     std_logic;
    iob25           : in     std_logic;
    iob26           : in     std_logic;
    iob27           : in     std_logic;
    iob28           : in     std_logic;
    iob29           : in     std_logic;
    iob3            : in     std_logic;
    iob30           : in     std_logic;
    iob31           : in     std_logic;
    iob32           : in     std_logic;
    iob33           : in     std_logic;
    iob34           : in     std_logic;
    iob35           : in     std_logic;
    iob36           : in     std_logic;
    iob37           : in     std_logic;
    iob38           : in     std_logic;
    iob39           : in     std_logic;
    iob4            : in     std_logic;
    iob40           : in     std_logic;
    iob41           : in     std_logic;
    iob42           : in     std_logic;
    iob43           : in     std_logic;
    iob44           : in     std_logic;
    iob45           : in     std_logic;
    iob46           : in     std_logic;
    iob47           : in     std_logic;
    iob5            : in     std_logic;
    iob6            : in     std_logic;
    iob7            : in     std_logic;
    iob8            : in     std_logic;
    iob9            : in     std_logic;
    ir0             : out    std_logic;
    ir1             : out    std_logic;
    ir10            : out    std_logic;
    ir11            : out    std_logic;
    ir12            : out    std_logic;
    ir13            : out    std_logic;
    ir14            : out    std_logic;
    ir15            : out    std_logic;
    ir16            : out    std_logic;
    ir17            : out    std_logic;
    ir18            : out    std_logic;
    ir19            : out    std_logic;
    ir2             : out    std_logic;
    ir20            : out    std_logic;
    ir21            : out    std_logic;
    ir22            : out    std_logic;
    ir23            : out    std_logic;
    ir24            : out    std_logic;
    ir25            : out    std_logic;
    ir26            : out    std_logic;
    ir27            : out    std_logic;
    ir28            : out    std_logic;
    ir29            : out    std_logic;
    ir3             : out    std_logic;
    ir30            : out    std_logic;
    ir31            : out    std_logic;
    ir32            : out    std_logic;
    ir33            : out    std_logic;
    ir34            : out    std_logic;
    ir35            : out    std_logic;
    ir36            : out    std_logic;
    ir37            : out    std_logic;
    ir38            : out    std_logic;
    ir39            : out    std_logic;
    ir4             : out    std_logic;
    ir40            : out    std_logic;
    ir41            : out    std_logic;
    ir42            : out    std_logic;
    ir43            : out    std_logic;
    ir44            : out    std_logic;
    ir45            : out    std_logic;
    ir46            : out    std_logic;
    ir47            : out    std_logic;
    ir48            : out    std_logic;
    ir5             : out    std_logic;
    ir6             : out    std_logic;
    ir7             : out    std_logic;
    ir8             : out    std_logic;
    ir9             : out    std_logic
  );
end entity cadr_ireg;
