library ieee;
use ieee.std_logic_1164.all;

package unsorted is

  component ic_16dummy port(dummy : in std_logic); end component;

end;

package body unsorted is

end;
