library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_stat is
  port (
    hi1        : in  std_logic;
    clk5a      : in  std_logic;
    iwr12      : in  std_logic;
    iwr13      : in  std_logic;
    iwr14      : in  std_logic;
    iwr15      : in  std_logic;
    gnd        : in  std_logic;
    \-ldstat\  : in  std_logic;
    \-stc12\   : out std_logic;
    st15       : out std_logic;
    st14       : out std_logic;
    st13       : out std_logic;
    st12       : out std_logic;
    \-stc16\   : out std_logic;
    iwr16      : in  std_logic;
    iwr17      : in  std_logic;
    iwr18      : in  std_logic;
    iwr19      : in  std_logic;
    st19       : out std_logic;
    st18       : out std_logic;
    st17       : out std_logic;
    st16       : out std_logic;
    \-stc20\   : out std_logic;
    iwr20      : in  std_logic;
    iwr21      : in  std_logic;
    iwr22      : in  std_logic;
    iwr23      : in  std_logic;
    st23       : out std_logic;
    st22       : out std_logic;
    st21       : out std_logic;
    st20       : out std_logic;
    \-stc24\   : out std_logic;
    iwr24      : in  std_logic;
    iwr25      : in  std_logic;
    iwr26      : in  std_logic;
    iwr27      : in  std_logic;
    st27       : out std_logic;
    st26       : out std_logic;
    st25       : out std_logic;
    st24       : out std_logic;
    \-stc28\   : out std_logic;
    iwr28      : in  std_logic;
    iwr29      : in  std_logic;
    iwr30      : in  std_logic;
    iwr31      : in  std_logic;
    st31       : out std_logic;
    st30       : out std_logic;
    st29       : out std_logic;
    st28       : out std_logic;
    \-stc32\   : out std_logic;
    \-spy.sth\ : in  std_logic;
    spy8       : out std_logic;
    spy9       : out std_logic;
    spy10      : out std_logic;
    spy11      : out std_logic;
    spy12      : out std_logic;
    spy13      : out std_logic;
    spy14      : out std_logic;
    spy15      : out std_logic;
    spy0       : out std_logic;
    spy1       : out std_logic;
    spy2       : out std_logic;
    spy3       : out std_logic;
    spy4       : out std_logic;
    spy5       : out std_logic;
    spy6       : out std_logic;
    spy7       : out std_logic;
    \-spy.stl\ : in  std_logic;
    st11       : out std_logic;
    st10       : out std_logic;
    st9        : out std_logic;
    st8        : out std_logic;
    st7        : out std_logic;
    st6        : out std_logic;
    st5        : out std_logic;
    st4        : out std_logic;
    st3        : out std_logic;
    st2        : out std_logic;
    st1        : out std_logic;
    st0        : out std_logic;
    iwr0       : in  std_logic;
    iwr1       : in  std_logic;
    iwr2       : in  std_logic;
    iwr3       : in  std_logic;
    \-statbit\ : in  std_logic;
    \-stc4\    : out std_logic;
    iwr4       : in  std_logic;
    iwr5       : in  std_logic;
    iwr6       : in  std_logic;
    iwr7       : in  std_logic;
    \-stc8\    : out std_logic;
    iwr8       : in  std_logic;
    iwr9       : in  std_logic;
    iwr10      : in  std_logic;
    iwr11      : in  std_logic);
end;

architecture ttl of cadr4_stat is
begin
  stat_1b01 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr12, i1 => iwr13, i2 => iwr14, i3 => iwr15, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc12\, o3 => st15, o2 => st14, o1 => st13, o0 => st12, co_n => \-stc16\);
  stat_1b02 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr16, i1 => iwr17, i2 => iwr18, i3 => iwr19, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc16\, o3 => st19, o2 => st18, o1 => st17, o0 => st16, co_n => \-stc20\);
  stat_1b03 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr20, i1 => iwr21, i2 => iwr22, i3 => iwr23, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc20\, o3 => st23, o2 => st22, o1 => st21, o0 => st20, co_n => \-stc24\);
  stat_1b04 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr24, i1 => iwr25, i2 => iwr26, i3 => iwr27, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc24\, o3 => st27, o2 => st26, o1 => st25, o0 => st24, co_n => \-stc28\);
  stat_1b05 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr28, i1 => iwr29, i2 => iwr30, i3 => iwr31, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc28\, o3 => st31, o2 => st30, o1 => st29, o0 => st28, co_n => \-stc32\);
  stat_1b06 : sn74ls244 port map(aenb_n => \-spy.sth\, ain0 => st31, bout3 => spy8, ain1 => st30, bout2 => spy9, ain2 => st29, bout1 => spy10, ain3 => st28, bout0 => spy11, bin0 => st27, aout3 => spy12, bin1 => st26, aout2 => spy13, bin2 => st25, aout1 => spy14, bin3 => st24, aout0 => spy15, benb_n => \-spy.sth\);
  stat_1b07 : sn74ls244 port map(aenb_n => \-spy.sth\, ain0 => st23, bout3 => spy0, ain1 => st22, bout2 => spy1, ain2 => st21, bout1 => spy2, ain3 => st20, bout0 => spy3, bin0 => st19, aout3 => spy4, bin1 => st18, aout2 => spy5, bin2 => st17, aout1 => spy6, bin3 => st16, aout0 => spy7, benb_n => \-spy.sth\);
  stat_1b08 : sn74ls244 port map(aenb_n => \-spy.stl\, ain0 => st15, bout3 => spy8, ain1 => st14, bout2 => spy9, ain2 => st13, bout1 => spy10, ain3 => st12, bout0 => spy11, bin0 => st11, aout3 => spy12, bin1 => st10, aout2 => spy13, bin2 => st9, aout1 => spy14, bin3 => st8, aout0 => spy15, benb_n => \-spy.stl\);
  stat_1b09 : sn74ls244 port map(aenb_n => \-spy.stl\, ain0 => st7, bout3 => spy0, ain1 => st6, bout2 => spy1, ain2 => st5, bout1 => spy2, ain3 => st4, bout0 => spy3, bin0 => st3, aout3 => spy4, bin1 => st2, aout2 => spy5, bin2 => st1, aout1 => spy6, bin3 => st0, aout0 => spy7, benb_n => \-spy.stl\);
  stat_1c03 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr0, i1 => iwr1, i2 => iwr2, i3 => iwr3, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-statbit\, o3 => st3, o2 => st2, o1 => st1, o0 => st0, co_n => \-stc4\);
  stat_1c04 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr4, i1 => iwr5, i2 => iwr6, i3 => iwr7, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc4\, o3 => st7, o2 => st6, o1 => st5, o0 => st4, co_n => \-stc8\);
  stat_1c05 : sn74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr8, i1 => iwr9, i2 => iwr10, i3 => iwr11, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc8\, o3 => st11, o2 => st10, o1 => st9, o0 => st8, co_n => \-stc12\);
end architecture;
