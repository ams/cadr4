library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sn7414 is
  port (
    g1a   : in  std_logic;
    g1q_n : out std_logic;
    g2a   : in  std_logic;
    g2q_n : out std_logic;
    g3a   : in  std_logic;
    g3q_n : out std_logic;
    g4q   : out std_logic;
    g4a   : in  std_logic;
    g5q_n : out std_logic;
    g5a   : in  std_logic;
    g6q_n : out std_logic;
    g6a   : in  std_logic
    );
end;

architecture ttl of sn7414 is
begin

end;
