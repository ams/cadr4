library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_9348 is
  port (
    i0  : in  std_logic;
    i1  : in  std_logic;
    i2  : in  std_logic;
    i3  : in  std_logic;
    i4  : in  std_logic;
    i5  : in  std_logic;
    i6  : in  std_logic;
    i7  : in  std_logic;
    i8  : in  std_logic;
    i9  : in  std_logic;
    i10 : in  std_logic;
    i11 : in  std_logic;
    pe  : out std_logic;
    po  : out std_logic
    );
end ic_9348;

architecture ttl of ic_9348 is
begin

end ttl;
