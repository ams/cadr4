library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn74260_tb is
end sn74260_tb;

architecture testbench of sn74260_tb is

begin

--  uut : sn74260 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
