-- CADR1_DIAG
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_diag is
  port (
    \-select spy\ : inout std_logic;
    \-spy read\ : out std_logic;
    \-spy write\ : out std_logic;
    \select spy\ : inout std_logic;
    \spy 0\ : inout std_logic;
    \spy 1\ : inout std_logic;
    \spy 10\ : inout std_logic;
    \spy 11\ : inout std_logic;
    \spy 12\ : inout std_logic;
    \spy 13\ : inout std_logic;
    \spy 14\ : inout std_logic;
    \spy 15\ : inout std_logic;
    \spy 2\ : inout std_logic;
    \spy 3\ : inout std_logic;
    \spy 4\ : inout std_logic;
    \spy 5\ : inout std_logic;
    \spy 6\ : inout std_logic;
    \spy 7\ : inout std_logic;
    \spy 8\ : inout std_logic;
    \spy 9\ : inout std_logic;
    \ub reg write pulse\ : in std_logic;
    ubrd : in std_logic;
    ubwr : inout std_logic;
    \udo 0\ : inout std_logic;
    \udo 1\ : inout std_logic;
    \udo 10\ : inout std_logic;
    \udo 11\ : inout std_logic;
    \udo 12\ : inout std_logic;
    \udo 13\ : inout std_logic;
    \udo 14\ : inout std_logic;
    \udo 15\ : inout std_logic;
    \udo 2\ : inout std_logic;
    \udo 3\ : inout std_logic;
    \udo 4\ : inout std_logic;
    \udo 5\ : inout std_logic;
    \udo 6\ : inout std_logic;
    \udo 7\ : inout std_logic;
    \udo 8\ : inout std_logic;
    \udo 9\ : inout std_logic
  );
end entity;
