library ieee;
use ieee.std_logic_1164.all;

entity icmem_iwrpar is
  port (
    iwr0            : in     std_logic;
    iwr1            : in     std_logic;
    iwr10           : in     std_logic;
    iwr11           : in     std_logic;
    iwr12           : in     std_logic;
    iwr13           : in     std_logic;
    iwr14           : in     std_logic;
    iwr15           : in     std_logic;
    iwr16           : in     std_logic;
    iwr17           : in     std_logic;
    iwr18           : in     std_logic;
    iwr19           : in     std_logic;
    iwr2            : in     std_logic;
    iwr20           : in     std_logic;
    iwr21           : in     std_logic;
    iwr22           : in     std_logic;
    iwr23           : in     std_logic;
    iwr24           : in     std_logic;
    iwr25           : in     std_logic;
    iwr26           : in     std_logic;
    iwr27           : in     std_logic;
    iwr28           : in     std_logic;
    iwr29           : in     std_logic;
    iwr3            : in     std_logic;
    iwr30           : in     std_logic;
    iwr31           : in     std_logic;
    iwr32           : in     std_logic;
    iwr33           : in     std_logic;
    iwr34           : in     std_logic;
    iwr35           : in     std_logic;
    iwr36           : in     std_logic;
    iwr37           : in     std_logic;
    iwr38           : in     std_logic;
    iwr39           : in     std_logic;
    iwr4            : in     std_logic;
    iwr40           : in     std_logic;
    iwr41           : in     std_logic;
    iwr42           : in     std_logic;
    iwr43           : in     std_logic;
    iwr44           : in     std_logic;
    iwr45           : in     std_logic;
    iwr46           : in     std_logic;
    iwr47           : in     std_logic;
    iwr5            : in     std_logic;
    iwr6            : in     std_logic;
    iwr7            : in     std_logic;
    iwr8            : in     std_logic;
    iwr9            : in     std_logic;
    iwr48           : out    std_logic;
    iwrp1           : out    std_logic;
    iwrp2           : out    std_logic;
    iwrp3           : out    std_logic;
    iwrp4           : out    std_logic
  );
end entity icmem_iwrpar;
