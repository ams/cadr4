library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_74260 is
  port (
    i1 : in  std_logic;
    i2 : in  std_logic;
    i3 : in  std_logic;
    o1 : out std_logic;
    i4 : in  std_logic;
    i5 : in  std_logic
    );
end ic_74260;

architecture ttl of ic_74260 is
begin

end ttl;
