library ieee;
use ieee.std_logic_1164.all;

entity helper_required_signals is
  port (
    \-halt\: out std_logic := '1';
    \-boot1\: out std_logic := '1'
  );
end entity;

architecture structural of helper_required_signals is
begin
end architecture;