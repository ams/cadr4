library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sip220_330_8 is
  port (
    r2 : in std_logic; -- 2
    r3 : in std_logic; -- 3
    r4 : in std_logic; -- 4
    r5 : in std_logic; -- 5
    r6 : in std_logic; -- 6
    r7 : in std_logic  -- 7
    );
end;

architecture ttl of sip220_330_8 is
begin
end;
