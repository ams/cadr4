library ieee;
use ieee.std_logic_1164.all;

entity cadr1_xapar is
  port (
    xao0            : in     std_logic;
    xao1            : in     std_logic;
    xao10           : in     std_logic;
    xao11           : in     std_logic;
    xao12           : in     std_logic;
    xao13           : in     std_logic;
    xao14           : in     std_logic;
    xao15           : in     std_logic;
    xao16           : in     std_logic;
    xao17           : in     std_logic;
    xao18           : in     std_logic;
    xao19           : in     std_logic;
    xao2            : in     std_logic;
    xao20           : in     std_logic;
    xao21           : in     std_logic;
    xao3            : in     std_logic;
    xao4            : in     std_logic;
    xao5            : in     std_logic;
    xao6            : in     std_logic;
    xao7            : in     std_logic;
    xao8            : in     std_logic;
    xao9            : in     std_logic;
    \xao par even\  : out    std_logic;
    \xao par odd\   : out    std_logic
  );
end entity cadr1_xapar;
