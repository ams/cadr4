library ieee;
use ieee.std_logic_1164.all;

entity cadr_amem0 is
  port (
    \-aadr0b\       : in     std_logic;
    \-aadr1b\       : in     std_logic;
    \-aadr2b\       : in     std_logic;
    \-aadr3b\       : in     std_logic;
    \-aadr4b\       : in     std_logic;
    \-aadr5b\       : in     std_logic;
    \-aadr6b\       : in     std_logic;
    \-aadr7b\       : in     std_logic;
    \-aadr8b\       : in     std_logic;
    \-aadr9b\       : in     std_logic;
    \-awpa\         : in     std_logic;
    \-awpb\         : in     std_logic;
    l16             : in     std_logic;
    l17             : in     std_logic;
    l18             : in     std_logic;
    l19             : in     std_logic;
    l20             : in     std_logic;
    l21             : in     std_logic;
    l22             : in     std_logic;
    l23             : in     std_logic;
    l24             : in     std_logic;
    l25             : in     std_logic;
    l26             : in     std_logic;
    l27             : in     std_logic;
    l28             : in     std_logic;
    l29             : in     std_logic;
    l30             : in     std_logic;
    l31             : in     std_logic;
    lparity         : in     std_logic;
    amem16          : out    std_logic;
    amem17          : out    std_logic;
    amem18          : out    std_logic;
    amem19          : out    std_logic;
    amem20          : out    std_logic;
    amem21          : out    std_logic;
    amem22          : out    std_logic;
    amem23          : out    std_logic;
    amem24          : out    std_logic;
    amem25          : out    std_logic;
    amem26          : out    std_logic;
    amem27          : out    std_logic;
    amem28          : out    std_logic;
    amem29          : out    std_logic;
    amem30          : out    std_logic;
    amem31          : out    std_logic;
    amemparity      : out    std_logic
  );
end entity;
