-- CADR1_UBD
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_ubd is
  port (
    \-ubd0\ : inout std_logic;
    \-ubd1\ : inout std_logic;
    \-ubd10\ : inout std_logic;
    \-ubd11\ : inout std_logic;
    \-ubd12\ : inout std_logic;
    \-ubd13\ : inout std_logic;
    \-ubd14\ : inout std_logic;
    \-ubd15\ : inout std_logic;
    \-ubd2\ : inout std_logic;
    \-ubd3\ : inout std_logic;
    \-ubd4\ : inout std_logic;
    \-ubd5\ : inout std_logic;
    \-ubd6\ : inout std_logic;
    \-ubd7\ : inout std_logic;
    \-ubd8\ : inout std_logic;
    \-ubd9\ : inout std_logic;
    \-ubdrive\ : inout std_logic;
    \-udi _ udo\ : in std_logic;
    \udi 0\ : in std_logic;
    \udi 1\ : in std_logic;
    \udi 10\ : in std_logic;
    \udi 11\ : in std_logic;
    \udi 12\ : in std_logic;
    \udi 13\ : in std_logic;
    \udi 14\ : in std_logic;
    \udi 15\ : in std_logic;
    \udi 2\ : in std_logic;
    \udi 3\ : in std_logic;
    \udi 4\ : in std_logic;
    \udi 5\ : in std_logic;
    \udi 6\ : in std_logic;
    \udi 7\ : in std_logic;
    \udi 8\ : in std_logic;
    \udi 9\ : in std_logic;
    udi0 : inout std_logic;
    udi1 : inout std_logic;
    udi10 : inout std_logic;
    udi11 : inout std_logic;
    udi12 : inout std_logic;
    udi13 : inout std_logic;
    udi14 : inout std_logic;
    udi15 : inout std_logic;
    udi2 : inout std_logic;
    udi3 : inout std_logic;
    udi4 : inout std_logic;
    udi5 : inout std_logic;
    udi6 : inout std_logic;
    udi7 : inout std_logic;
    udi8 : inout std_logic;
    udi9 : inout std_logic;
    \udo 0\ : out std_logic;
    \udo 1\ : out std_logic;
    \udo 10\ : out std_logic;
    \udo 11\ : out std_logic;
    \udo 12\ : out std_logic;
    \udo 13\ : out std_logic;
    \udo 14\ : out std_logic;
    \udo 15\ : out std_logic;
    \udo 2\ : out std_logic;
    \udo 3\ : out std_logic;
    \udo 4\ : out std_logic;
    \udo 5\ : out std_logic;
    \udo 6\ : out std_logic;
    \udo 7\ : out std_logic;
    \udo 8\ : out std_logic;
    \udo 9\ : out std_logic;
    udo0 : inout std_logic;
    udo1 : inout std_logic;
    udo10 : inout std_logic;
    udo11 : inout std_logic;
    udo12 : inout std_logic;
    udo13 : inout std_logic;
    udo14 : inout std_logic;
    udo15 : inout std_logic;
    udo2 : inout std_logic;
    udo3 : inout std_logic;
    udo4 : inout std_logic;
    udo5 : inout std_logic;
    udo6 : inout std_logic;
    udo7 : inout std_logic;
    udo8 : inout std_logic;
    udo9 : inout std_logic
  );
end entity;
