-- The MIT CADR

library ieee;
use ieee.std_logic_1164.all;

use std.env.finish;

use work.cadr_book.all;
use work.icmem_book.all;

entity cadr_tb is
end;

architecture structural of cadr_tb is
  signal \-a31\ : std_logic := '0';
  signal \-aadr0a\ : std_logic := '0';
  signal \-aadr0b\ : std_logic := '0';
  signal \-aadr1a\ : std_logic := '0';
  signal \-aadr1b\ : std_logic := '0';
  signal \-aadr2a\ : std_logic := '0';
  signal \-aadr2b\ : std_logic := '0';
  signal \-aadr3a\ : std_logic := '0';
  signal \-aadr3b\ : std_logic := '0';
  signal \-aadr4a\ : std_logic := '0';
  signal \-aadr4b\ : std_logic := '0';
  signal \-aadr5a\ : std_logic := '0';
  signal \-aadr5b\ : std_logic := '0';
  signal \-aadr6a\ : std_logic := '0';
  signal \-aadr6b\ : std_logic := '0';
  signal \-aadr7a\ : std_logic := '0';
  signal \-aadr7b\ : std_logic := '0';
  signal \-aadr8a\ : std_logic := '0';
  signal \-aadr8b\ : std_logic := '0';
  signal \-aadr9a\ : std_logic := '0';
  signal \-aadr9b\ : std_logic := '0';
  signal \-adrpar\ : std_logic := '0';
  signal \-alu31\ : std_logic := '0';
  signal \-alu32\ : std_logic := '0';
  signal \-aluf0\ : std_logic := '0';
  signal \-aluf1\ : std_logic := '0';
  signal \-aluf2\ : std_logic := '0';
  signal \-aluf3\ : std_logic := '0';
  signal \-alumode\ : std_logic := '0';
  signal \-amemenb\ : std_logic := '0';
  signal \-apass\ : std_logic := '0';
  signal \-apassenb\ : std_logic := '0';
  signal \-ape\ : std_logic := '0';
  signal \-awpa\ : std_logic := '0';
  signal \-awpb\ : std_logic := '0';
  signal \-awpc\ : std_logic := '0';
  signal \-boot1\ : std_logic := '0';
  signal \-boot2\ : std_logic := '0';
  signal \-boot\ : std_logic := '0';
  signal \-bus.reset\ : std_logic := '0';
  signal \-busint.lm.reset\ : std_logic := '0';
  signal \-cin0\ : std_logic := '0';
  signal \-cin12\ : std_logic := '0';
  signal \-cin16\ : std_logic := '0';
  signal \-cin20\ : std_logic := '0';
  signal \-cin24\ : std_logic := '0';
  signal \-cin28\ : std_logic := '0';
  signal \-cin32\ : std_logic := '0';
  signal \-cin4\ : std_logic := '0';
  signal \-cin8\ : std_logic := '0';
  signal \-clk0\ : std_logic := '0';
  signal \-clk1\ : std_logic := '0';
  signal \-clk2a\ : std_logic := '0';
  signal \-clk2c\ : std_logic := '0';
  signal \-clk3a\ : std_logic := '0';
  signal \-clk3d\ : std_logic := '0';
  signal \-clk3g\ : std_logic := '0';
  signal \-clk4a\ : std_logic := '0';
  signal \-clk4d\ : std_logic := '0';
  signal \-clk4e\ : std_logic := '0';
  signal \-clk5\ : std_logic := '0';
  signal \-clock_reset_a\ : std_logic := '0';
  signal \-clock_reset_b\ : std_logic := '0';
  signal \-dadr0a\ : std_logic := '0';
  signal \-dadr0b\ : std_logic := '0';
  signal \-dadr0c\ : std_logic := '0';
  signal \-dadr10a\ : std_logic := '0';
  signal \-dadr10c\ : std_logic := '0';
  signal \-dadr1a\ : std_logic := '0';
  signal \-dadr1b\ : std_logic := '0';
  signal \-dadr1c\ : std_logic := '0';
  signal \-dadr2a\ : std_logic := '0';
  signal \-dadr2b\ : std_logic := '0';
  signal \-dadr2c\ : std_logic := '0';
  signal \-dadr3a\ : std_logic := '0';
  signal \-dadr3b\ : std_logic := '0';
  signal \-dadr3c\ : std_logic := '0';
  signal \-dadr4a\ : std_logic := '0';
  signal \-dadr4b\ : std_logic := '0';
  signal \-dadr4c\ : std_logic := '0';
  signal \-dadr5a\ : std_logic := '0';
  signal \-dadr5b\ : std_logic := '0';
  signal \-dadr5c\ : std_logic := '0';
  signal \-dadr6a\ : std_logic := '0';
  signal \-dadr6b\ : std_logic := '0';
  signal \-dadr6c\ : std_logic := '0';
  signal \-dadr7a\ : std_logic := '0';
  signal \-dadr7b\ : std_logic := '0';
  signal \-dadr7c\ : std_logic := '0';
  signal \-dadr8a\ : std_logic := '0';
  signal \-dadr8b\ : std_logic := '0';
  signal \-dadr8c\ : std_logic := '0';
  signal \-dadr9a\ : std_logic := '0';
  signal \-dadr9b\ : std_logic := '0';
  signal \-dadr9c\ : std_logic := '0';
  signal \-dbread\ : std_logic := '0';
  signal \-dbwrite\ : std_logic := '0';
  signal \-destimod0\ : std_logic := '0';
  signal \-destimod1\ : std_logic := '0';
  signal \-destintctl\ : std_logic := '0';
  signal \-destlc\ : std_logic := '0';
  signal \-destmdr\ : std_logic := '0';
  signal \-destmem\ : std_logic := '0';
  signal \-destpdl(p)\ : std_logic := '0';
  signal \-destpdl(x)\ : std_logic := '0';
  signal \-destpdlp\ : std_logic := '0';
  signal \-destpdltop\ : std_logic := '0';
  signal \-destpdlx\ : std_logic := '0';
  signal \-destspc\ : std_logic := '0';
  signal \-destspcd\ : std_logic := '0';
  signal \-destvma\ : std_logic := '0';
  signal \-dfall\ : std_logic := '0';
  signal \-div\ : std_logic := '0';
  signal \-divposlasttime\ : std_logic := '0';
  signal \-dmapbenb\ : std_logic := '0';
  signal \-dp\ : std_logic := '0';
  signal \-dparh\ : std_logic := '0';
  signal \-dpe\ : std_logic := '0';
  signal \-dr\ : std_logic := '0';
  signal \-dwea\ : std_logic := '0';
  signal \-dweb\ : std_logic := '0';
  signal \-dwec\ : std_logic := '0';
  signal \-errhalt\ : std_logic := '0';
  signal \-funct0\ : std_logic := '0';
  signal \-funct1\ : std_logic := '0';
  signal \-funct2\ : std_logic := '0';
  signal \-funct3\ : std_logic := '0';
  signal \-halt\ : std_logic := '0';
  signal \-halted\ : std_logic := '0';
  signal \-hang\ : std_logic := '0';
  signal \-higherr\ : std_logic := '0';
  signal \-ice0a\ : std_logic := '0';
  signal \-ice0b\ : std_logic := '0';
  signal \-ice0c\ : std_logic := '0';
  signal \-ice0d\ : std_logic := '0';
  signal \-ice1a\ : std_logic := '0';
  signal \-ice1b\ : std_logic := '0';
  signal \-ice1c\ : std_logic := '0';
  signal \-ice1d\ : std_logic := '0';
  signal \-ice2a\ : std_logic := '0';
  signal \-ice2b\ : std_logic := '0';
  signal \-ice2c\ : std_logic := '0';
  signal \-ice2d\ : std_logic := '0';
  signal \-ice3a\ : std_logic := '0';
  signal \-ice3b\ : std_logic := '0';
  signal \-ice3c\ : std_logic := '0';
  signal \-ice3d\ : std_logic := '0';
  signal \-idebug\ : std_logic := '0';
  signal \-ifetch\ : std_logic := '0';
  signal \-ignpar\ : std_logic := '0';
  signal \-ignpopj\ : std_logic := '0';
  signal \-ilong\ : std_logic := '0';
  signal \-imodd\ : std_logic := '0';
  signal \-inop\ : std_logic := '0';
  signal \-ipe\ : std_logic := '0';
  signal \-ipopj\ : std_logic := '0';
  signal \-ir0\ : std_logic := '0';
  signal \-ir12\ : std_logic := '0';
  signal \-ir13\ : std_logic := '0';
  signal \-ir1\ : std_logic := '0';
  signal \-ir22\ : std_logic := '0';
  signal \-ir25\ : std_logic := '0';
  signal \-ir2\ : std_logic := '0';
  signal \-ir31\ : std_logic := '0';
  signal \-ir3\ : std_logic := '0';
  signal \-ir4\ : std_logic := '0';
  signal \-ir6\ : std_logic := '0';
  signal \-ir8\ : std_logic := '0';
  signal \-iralu\ : std_logic := '0';
  signal \-irbyte\ : std_logic := '0';
  signal \-irdisp\ : std_logic := '0';
  signal \-irjump\ : std_logic := '0';
  signal \-iwea\ : std_logic := '0';
  signal \-iweb\ : std_logic := '0';
  signal \-iwec\ : std_logic := '0';
  signal \-iwed\ : std_logic := '0';
  signal \-iwee\ : std_logic := '0';
  signal \-iwef\ : std_logic := '0';
  signal \-iweg\ : std_logic := '0';
  signal \-iweh\ : std_logic := '0';
  signal \-iwei\ : std_logic := '0';
  signal \-iwej\ : std_logic := '0';
  signal \-iwek\ : std_logic := '0';
  signal \-iwel\ : std_logic := '0';
  signal \-iwem\ : std_logic := '0';
  signal \-iwen\ : std_logic := '0';
  signal \-iweo\ : std_logic := '0';
  signal \-iwep\ : std_logic := '0';
  signal \-iwrited\ : std_logic := '0';
  signal \-iwriteda\ : std_logic := '0';
  signal \-jcond\ : std_logic := '0';
  signal \-lc_modifies_mrot\ : std_logic := '0';
  signal \-lcdrive\ : std_logic := '0';
  signal \-lcinc\ : std_logic := '0';
  signal \-lcry11\ : std_logic := '0';
  signal \-lcry15\ : std_logic := '0';
  signal \-lcry19\ : std_logic := '0';
  signal \-lcry23\ : std_logic := '0';
  signal \-lcry3\ : std_logic := '0';
  signal \-lcry7\ : std_logic := '0';
  signal \-ldclk\ : std_logic := '0';
  signal \-lddbirh\ : std_logic := '0';
  signal \-lddbirl\ : std_logic := '0';
  signal \-lddbirm\ : std_logic := '0';
  signal \-ldmode\ : std_logic := '0';
  signal \-ldopc\ : std_logic := '0';
  signal \-ldstat\ : std_logic := '0';
  signal \-loadmd\ : std_logic := '0';
  signal \-lowerhighok\ : std_logic := '0';
  signal \-lparity\ : std_logic := '0';
  signal \-lparm\ : std_logic := '0';
  signal \-lpc.hold\ : std_logic := '0';
  signal \-lvmo22\ : std_logic := '0';
  signal \-lvmo23\ : std_logic := '0';
  signal \-machrun\ : std_logic := '0';
  signal \-machruna\ : std_logic := '0';
  signal \-madr0a\ : std_logic := '0';
  signal \-madr0b\ : std_logic := '0';
  signal \-madr1a\ : std_logic := '0';
  signal \-madr1b\ : std_logic := '0';
  signal \-madr2a\ : std_logic := '0';
  signal \-madr2b\ : std_logic := '0';
  signal \-madr3a\ : std_logic := '0';
  signal \-madr3b\ : std_logic := '0';
  signal \-madr4a\ : std_logic := '0';
  signal \-madr4b\ : std_logic := '0';
  signal \-mapdrive\ : std_logic := '0';
  signal \-mapi10a\ : std_logic := '0';
  signal \-mapi10b\ : std_logic := '0';
  signal \-mapi11a\ : std_logic := '0';
  signal \-mapi11b\ : std_logic := '0';
  signal \-mapi12a\ : std_logic := '0';
  signal \-mapi12b\ : std_logic := '0';
  signal \-mapi23\ : std_logic := '0';
  signal \-mapi8a\ : std_logic := '0';
  signal \-mapi8b\ : std_logic := '0';
  signal \-mapi9a\ : std_logic := '0';
  signal \-mapi9b\ : std_logic := '0';
  signal \-mbusy.sync\ : std_logic := '0';
  signal \-mclk0\ : std_logic := '0';
  signal \-mclk1\ : std_logic := '0';
  signal \-mclk5\ : std_logic := '0';
  signal \-md0\ : std_logic := '0';
  signal \-md10\ : std_logic := '0';
  signal \-md11\ : std_logic := '0';
  signal \-md12\ : std_logic := '0';
  signal \-md13\ : std_logic := '0';
  signal \-md14\ : std_logic := '0';
  signal \-md15\ : std_logic := '0';
  signal \-md16\ : std_logic := '0';
  signal \-md17\ : std_logic := '0';
  signal \-md18\ : std_logic := '0';
  signal \-md19\ : std_logic := '0';
  signal \-md1\ : std_logic := '0';
  signal \-md20\ : std_logic := '0';
  signal \-md21\ : std_logic := '0';
  signal \-md22\ : std_logic := '0';
  signal \-md23\ : std_logic := '0';
  signal \-md24\ : std_logic := '0';
  signal \-md25\ : std_logic := '0';
  signal \-md26\ : std_logic := '0';
  signal \-md27\ : std_logic := '0';
  signal \-md28\ : std_logic := '0';
  signal \-md29\ : std_logic := '0';
  signal \-md2\ : std_logic := '0';
  signal \-md30\ : std_logic := '0';
  signal \-md31\ : std_logic := '0';
  signal \-md3\ : std_logic := '0';
  signal \-md4\ : std_logic := '0';
  signal \-md5\ : std_logic := '0';
  signal \-md6\ : std_logic := '0';
  signal \-md7\ : std_logic := '0';
  signal \-md8\ : std_logic := '0';
  signal \-md9\ : std_logic := '0';
  signal \-mddrive\ : std_logic := '0';
  signal \-mds0\ : std_logic := '0';
  signal \-mds10\ : std_logic := '0';
  signal \-mds11\ : std_logic := '0';
  signal \-mds12\ : std_logic := '0';
  signal \-mds13\ : std_logic := '0';
  signal \-mds14\ : std_logic := '0';
  signal \-mds15\ : std_logic := '0';
  signal \-mds16\ : std_logic := '0';
  signal \-mds17\ : std_logic := '0';
  signal \-mds18\ : std_logic := '0';
  signal \-mds19\ : std_logic := '0';
  signal \-mds1\ : std_logic := '0';
  signal \-mds20\ : std_logic := '0';
  signal \-mds21\ : std_logic := '0';
  signal \-mds22\ : std_logic := '0';
  signal \-mds23\ : std_logic := '0';
  signal \-mds24\ : std_logic := '0';
  signal \-mds25\ : std_logic := '0';
  signal \-mds26\ : std_logic := '0';
  signal \-mds27\ : std_logic := '0';
  signal \-mds28\ : std_logic := '0';
  signal \-mds29\ : std_logic := '0';
  signal \-mds2\ : std_logic := '0';
  signal \-mds30\ : std_logic := '0';
  signal \-mds31\ : std_logic := '0';
  signal \-mds3\ : std_logic := '0';
  signal \-mds4\ : std_logic := '0';
  signal \-mds5\ : std_logic := '0';
  signal \-mds6\ : std_logic := '0';
  signal \-mds7\ : std_logic := '0';
  signal \-mds8\ : std_logic := '0';
  signal \-mds9\ : std_logic := '0';
  signal \-memack\ : std_logic := '0';
  signal \-memdrive.a\ : std_logic := '0';
  signal \-memdrive.b\ : std_logic := '0';
  signal \-memgrant\ : std_logic := '0';
  signal \-memop\ : std_logic := '0';
  signal \-memparok\ : std_logic := '0';
  signal \-mempe\ : std_logic := '0';
  signal \-memprepare\ : std_logic := '0';
  signal \-memrd\ : std_logic := '0';
  signal \-memrq\ : std_logic := '0';
  signal \-memstart\ : std_logic := '0';
  signal \-memwr\ : std_logic := '0';
  signal \-mfdrive\ : std_logic := '0';
  signal \-mfinish\ : std_logic := '0';
  signal \-mfinishd\ : std_logic := '0';
  signal \-mpass\ : std_logic := '0';
  signal \-mpassl\ : std_logic := '0';
  signal \-mpassm\ : std_logic := '0';
  signal \-mpe\ : std_logic := '0';
  signal \-mr\ : std_logic := '0';
  signal \-mul\ : std_logic := '0';
  signal \-mulnop\ : std_logic := '0';
  signal \-mwpa\ : std_logic := '0';
  signal \-mwpb\ : std_logic := '0';
  signal \-needfetch\ : std_logic := '0';
  signal \-newlc.in\ : std_logic := '0';
  signal \-newlc\ : std_logic := '0';
  signal \-nop11\ : std_logic := '0';
  signal \-nop\ : std_logic := '0';
  signal \-nopa\ : std_logic := '0';
  signal \-opcclk\ : std_logic := '0';
  signal \-opcdrive\ : std_logic := '0';
  signal \-opcinh\ : std_logic := '0';
  signal \-parerr\ : std_logic := '0';
  signal \-pc12b\ : std_logic := '0';
  signal \-pc13b\ : std_logic := '0';
  signal \-pcb0\ : std_logic := '0';
  signal \-pcb10\ : std_logic := '0';
  signal \-pcb11\ : std_logic := '0';
  signal \-pcb1\ : std_logic := '0';
  signal \-pcb2\ : std_logic := '0';
  signal \-pcb3\ : std_logic := '0';
  signal \-pcb4\ : std_logic := '0';
  signal \-pcb5\ : std_logic := '0';
  signal \-pcb6\ : std_logic := '0';
  signal \-pcb7\ : std_logic := '0';
  signal \-pcb8\ : std_logic := '0';
  signal \-pcb9\ : std_logic := '0';
  signal \-pcc0\ : std_logic := '0';
  signal \-pcc10\ : std_logic := '0';
  signal \-pcc11\ : std_logic := '0';
  signal \-pcc1\ : std_logic := '0';
  signal \-pcc2\ : std_logic := '0';
  signal \-pcc3\ : std_logic := '0';
  signal \-pcc4\ : std_logic := '0';
  signal \-pcc5\ : std_logic := '0';
  signal \-pcc6\ : std_logic := '0';
  signal \-pcc7\ : std_logic := '0';
  signal \-pcc8\ : std_logic := '0';
  signal \-pcc9\ : std_logic := '0';
  signal \-pdla0a\ : std_logic := '0';
  signal \-pdla0b\ : std_logic := '0';
  signal \-pdla1a\ : std_logic := '0';
  signal \-pdla1b\ : std_logic := '0';
  signal \-pdla2a\ : std_logic := '0';
  signal \-pdla2b\ : std_logic := '0';
  signal \-pdla3a\ : std_logic := '0';
  signal \-pdla3b\ : std_logic := '0';
  signal \-pdla4a\ : std_logic := '0';
  signal \-pdla4b\ : std_logic := '0';
  signal \-pdla5a\ : std_logic := '0';
  signal \-pdla5b\ : std_logic := '0';
  signal \-pdla6a\ : std_logic := '0';
  signal \-pdla6b\ : std_logic := '0';
  signal \-pdla7a\ : std_logic := '0';
  signal \-pdla7b\ : std_logic := '0';
  signal \-pdla8a\ : std_logic := '0';
  signal \-pdla8b\ : std_logic := '0';
  signal \-pdla9a\ : std_logic := '0';
  signal \-pdla9b\ : std_logic := '0';
  signal \-pdlcnt\ : std_logic := '0';
  signal \-pdlcry3\ : std_logic := '0';
  signal \-pdlcry7\ : std_logic := '0';
  signal \-pdldrive\ : std_logic := '0';
  signal \-pdlpa\ : std_logic := '0';
  signal \-pdlpb\ : std_logic := '0';
  signal \-pdlpe\ : std_logic := '0';
  signal \-pdlwrited\ : std_logic := '0';
  signal \-pfr\ : std_logic := '0';
  signal \-pfw\ : std_logic := '0';
  signal \-pma10\ : std_logic := '0';
  signal \-pma11\ : std_logic := '0';
  signal \-pma12\ : std_logic := '0';
  signal \-pma13\ : std_logic := '0';
  signal \-pma14\ : std_logic := '0';
  signal \-pma15\ : std_logic := '0';
  signal \-pma16\ : std_logic := '0';
  signal \-pma17\ : std_logic := '0';
  signal \-pma18\ : std_logic := '0';
  signal \-pma19\ : std_logic := '0';
  signal \-pma20\ : std_logic := '0';
  signal \-pma21\ : std_logic := '0';
  signal \-pma8\ : std_logic := '0';
  signal \-pma9\ : std_logic := '0';
  signal \-popj\ : std_logic := '0';
  signal \-power_reset\ : std_logic := '0';
  signal \-ppdrive\ : std_logic := '0';
  signal \-prog.reset\ : std_logic := '0';
  signal \-promce0\ : std_logic := '0';
  signal \-promce1\ : std_logic := '0';
  signal \-promdisabled\ : std_logic := '0';
  signal \-promenable\ : std_logic := '0';
  signal \-prompc0\ : std_logic := '0';
  signal \-prompc1\ : std_logic := '0';
  signal \-prompc2\ : std_logic := '0';
  signal \-prompc3\ : std_logic := '0';
  signal \-prompc4\ : std_logic := '0';
  signal \-prompc5\ : std_logic := '0';
  signal \-prompc6\ : std_logic := '0';
  signal \-prompc7\ : std_logic := '0';
  signal \-prompc8\ : std_logic := '0';
  signal \-prompc9\ : std_logic := '0';
  signal \-pwidx\ : std_logic := '0';
  signal \-pwpa\ : std_logic := '0';
  signal \-pwpb\ : std_logic := '0';
  signal \-pwpc\ : std_logic := '0';
  signal \-qdrive\ : std_logic := '0';
  signal \-rdfinish\ : std_logic := '0';
  signal \-reset\ : std_logic := '0';
  signal \-run\ : std_logic := '0';
  signal \-s4\ : std_logic := '0';
  signal \-sh3\ : std_logic := '0';
  signal \-sh4\ : std_logic := '0';
  signal \-spccry\ : std_logic := '0';
  signal \-spcdrive\ : std_logic := '0';
  signal \-spcnt\ : std_logic := '0';
  signal \-spcpass\ : std_logic := '0';
  signal \-spcwparl\ : std_logic := '0';
  signal \-spcwpass\ : std_logic := '0';
  signal \-spe\ : std_logic := '0';
  signal \-specalu\ : std_logic := '0';
  signal \-spop\ : std_logic := '0';
  signal \-spush\ : std_logic := '0';
  signal \-spushd\ : std_logic := '0';
  signal \-spy.ah\ : std_logic := '0';
  signal \-spy.al\ : std_logic := '0';
  signal \-spy.flag1\ : std_logic := '0';
  signal \-spy.flag2\ : std_logic := '0';
  signal \-spy.irh\ : std_logic := '0';
  signal \-spy.irl\ : std_logic := '0';
  signal \-spy.irm\ : std_logic := '0';
  signal \-spy.mh\ : std_logic := '0';
  signal \-spy.ml\ : std_logic := '0';
  signal \-spy.obh\ : std_logic := '0';
  signal \-spy.obl\ : std_logic := '0';
  signal \-spy.opc\ : std_logic := '0';
  signal \-spy.pc\ : std_logic := '0';
  signal \-spy.sth\ : std_logic := '0';
  signal \-spy.stl\ : std_logic := '0';
  signal \-sr\ : std_logic := '0';
  signal \-srcdc\ : std_logic := '0';
  signal \-srclc\ : std_logic := '0';
  signal \-srcm\ : std_logic := '0';
  signal \-srcmap\ : std_logic := '0';
  signal \-srcmd\ : std_logic := '0';
  signal \-srcopc\ : std_logic := '0';
  signal \-srcpdlidx\ : std_logic := '0';
  signal \-srcpdlpop\ : std_logic := '0';
  signal \-srcpdlptr\ : std_logic := '0';
  signal \-srcpdltop\ : std_logic := '0';
  signal \-srcq\ : std_logic := '0';
  signal \-srcspc\ : std_logic := '0';
  signal \-srcspcpop\ : std_logic := '0';
  signal \-srcspcpopreal\ : std_logic := '0';
  signal \-srcvma\ : std_logic := '0';
  signal \-ssdone\ : std_logic := '0';
  signal \-statbit\ : std_logic := '0';
  signal \-stathalt\ : std_logic := '0';
  signal \-stc12\ : std_logic := '0';
  signal \-stc16\ : std_logic := '0';
  signal \-stc20\ : std_logic := '0';
  signal \-stc24\ : std_logic := '0';
  signal \-stc28\ : std_logic := '0';
  signal \-stc32\ : std_logic := '0';
  signal \-stc4\ : std_logic := '0';
  signal \-stc8\ : std_logic := '0';
  signal \-step\ : std_logic := '0';
  signal \-swpa\ : std_logic := '0';
  signal \-swpb\ : std_logic := '0';
  signal \-tpclk\ : std_logic := '0';
  signal \-tpdone\ : std_logic := '0';
  signal \-tpr0\ : std_logic := '0';
  signal \-tpr100\ : std_logic := '0';
  signal \-tpr105\ : std_logic := '0';
  signal \-tpr10\ : std_logic := '0';
  signal \-tpr110\ : std_logic := '0';
  signal \-tpr115\ : std_logic := '0';
  signal \-tpr120\ : std_logic := '0';
  signal \-tpr120a\ : std_logic := '0';
  signal \-tpr125\ : std_logic := '0';
  signal \-tpr140\ : std_logic := '0';
  signal \-tpr15\ : std_logic := '0';
  signal \-tpr160\ : std_logic := '0';
  signal \-tpr180\ : std_logic := '0';
  signal \-tpr200\ : std_logic := '0';
  signal \-tpr20\ : std_logic := '0';
  signal \-tpr20a\ : std_logic := '0';
  signal \-tpr25\ : std_logic := '0';
  signal \-tpr40\ : std_logic := '0';
  signal \-tpr5\ : std_logic := '0';
  signal \-tpr60\ : std_logic := '0';
  signal \-tpr65\ : std_logic := '0';
  signal \-tpr70\ : std_logic := '0';
  signal \-tpr75\ : std_logic := '0';
  signal \-tpr80\ : std_logic := '0';
  signal \-tpr80a\ : std_logic := '0';
  signal \-tpr85\ : std_logic := '0';
  signal \-tprend\ : std_logic := '0';
  signal \-tptse\ : std_logic := '0';
  signal \-tpw10\ : std_logic := '0';
  signal \-tpw20\ : std_logic := '0';
  signal \-tpw25\ : std_logic := '0';
  signal \-tpw30\ : std_logic := '0';
  signal \-tpw30a\ : std_logic := '0';
  signal \-tpw35\ : std_logic := '0';
  signal \-tpw40\ : std_logic := '0';
  signal \-tpw40a\ : std_logic := '0';
  signal \-tpw45\ : std_logic := '0';
  signal \-tpw50\ : std_logic := '0';
  signal \-tpw55\ : std_logic := '0';
  signal \-tpw60\ : std_logic := '0';
  signal \-tpw65\ : std_logic := '0';
  signal \-tpw70\ : std_logic := '0';
  signal \-tpw75\ : std_logic := '0';
  signal \-trap\ : std_logic := '0';
  signal \-trapenb\ : std_logic := '0';
  signal \-tse1\ : std_logic := '0';
  signal \-tse2\ : std_logic := '0';
  signal \-tse3\ : std_logic := '0';
  signal \-tse4\ : std_logic := '0';
  signal \-upperhighok\ : std_logic := '0';
  signal \-use.map\ : std_logic := '0';
  signal \-v0pe\ : std_logic := '0';
  signal \-v1pe\ : std_logic := '0';
  signal \-vm0wpa\ : std_logic := '0';
  signal \-vm0wpb\ : std_logic := '0';
  signal \-vm1lpar\ : std_logic := '0';
  signal \-vm1wpa\ : std_logic := '0';
  signal \-vm1wpb\ : std_logic := '0';
  signal \-vma0\ : std_logic := '0';
  signal \-vma10\ : std_logic := '0';
  signal \-vma11\ : std_logic := '0';
  signal \-vma12\ : std_logic := '0';
  signal \-vma13\ : std_logic := '0';
  signal \-vma14\ : std_logic := '0';
  signal \-vma15\ : std_logic := '0';
  signal \-vma16\ : std_logic := '0';
  signal \-vma17\ : std_logic := '0';
  signal \-vma18\ : std_logic := '0';
  signal \-vma19\ : std_logic := '0';
  signal \-vma1\ : std_logic := '0';
  signal \-vma20\ : std_logic := '0';
  signal \-vma21\ : std_logic := '0';
  signal \-vma22\ : std_logic := '0';
  signal \-vma23\ : std_logic := '0';
  signal \-vma24\ : std_logic := '0';
  signal \-vma25\ : std_logic := '0';
  signal \-vma26\ : std_logic := '0';
  signal \-vma27\ : std_logic := '0';
  signal \-vma28\ : std_logic := '0';
  signal \-vma29\ : std_logic := '0';
  signal \-vma2\ : std_logic := '0';
  signal \-vma30\ : std_logic := '0';
  signal \-vma31\ : std_logic := '0';
  signal \-vma3\ : std_logic := '0';
  signal \-vma4\ : std_logic := '0';
  signal \-vma5\ : std_logic := '0';
  signal \-vma6\ : std_logic := '0';
  signal \-vma7\ : std_logic := '0';
  signal \-vma8\ : std_logic := '0';
  signal \-vma9\ : std_logic := '0';
  signal \-vmadrive\ : std_logic := '0';
  signal \-vmaenb\ : std_logic := '0';
  signal \-vmaok\ : std_logic := '0';
  signal \-vmap0\ : std_logic := '0';
  signal \-vmap1\ : std_logic := '0';
  signal \-vmap2\ : std_logic := '0';
  signal \-vmap3\ : std_logic := '0';
  signal \-vmap4\ : std_logic := '0';
  signal \-vmas0\ : std_logic := '0';
  signal \-vmas10\ : std_logic := '0';
  signal \-vmas11\ : std_logic := '0';
  signal \-vmas12\ : std_logic := '0';
  signal \-vmas13\ : std_logic := '0';
  signal \-vmas14\ : std_logic := '0';
  signal \-vmas15\ : std_logic := '0';
  signal \-vmas16\ : std_logic := '0';
  signal \-vmas17\ : std_logic := '0';
  signal \-vmas18\ : std_logic := '0';
  signal \-vmas19\ : std_logic := '0';
  signal \-vmas1\ : std_logic := '0';
  signal \-vmas20\ : std_logic := '0';
  signal \-vmas21\ : std_logic := '0';
  signal \-vmas22\ : std_logic := '0';
  signal \-vmas23\ : std_logic := '0';
  signal \-vmas24\ : std_logic := '0';
  signal \-vmas25\ : std_logic := '0';
  signal \-vmas26\ : std_logic := '0';
  signal \-vmas27\ : std_logic := '0';
  signal \-vmas28\ : std_logic := '0';
  signal \-vmas29\ : std_logic := '0';
  signal \-vmas2\ : std_logic := '0';
  signal \-vmas30\ : std_logic := '0';
  signal \-vmas31\ : std_logic := '0';
  signal \-vmas3\ : std_logic := '0';
  signal \-vmas4\ : std_logic := '0';
  signal \-vmas5\ : std_logic := '0';
  signal \-vmas6\ : std_logic := '0';
  signal \-vmas7\ : std_logic := '0';
  signal \-vmas8\ : std_logic := '0';
  signal \-vmas9\ : std_logic := '0';
  signal \-vmo0\ : std_logic := '0';
  signal \-vmo10\ : std_logic := '0';
  signal \-vmo11\ : std_logic := '0';
  signal \-vmo12\ : std_logic := '0';
  signal \-vmo13\ : std_logic := '0';
  signal \-vmo14\ : std_logic := '0';
  signal \-vmo15\ : std_logic := '0';
  signal \-vmo16\ : std_logic := '0';
  signal \-vmo17\ : std_logic := '0';
  signal \-vmo18\ : std_logic := '0';
  signal \-vmo19\ : std_logic := '0';
  signal \-vmo1\ : std_logic := '0';
  signal \-vmo20\ : std_logic := '0';
  signal \-vmo21\ : std_logic := '0';
  signal \-vmo22\ : std_logic := '0';
  signal \-vmo23\ : std_logic := '0';
  signal \-vmo2\ : std_logic := '0';
  signal \-vmo3\ : std_logic := '0';
  signal \-vmo4\ : std_logic := '0';
  signal \-vmo5\ : std_logic := '0';
  signal \-vmo6\ : std_logic := '0';
  signal \-vmo7\ : std_logic := '0';
  signal \-vmo8\ : std_logic := '0';
  signal \-vmo9\ : std_logic := '0';
  signal \-wait\ : std_logic := '0';
  signal \-wmap\ : std_logic := '0';
  signal \-wmapd\ : std_logic := '0';
  signal \-wp1\ : std_logic := '0';
  signal \-wp2\ : std_logic := '0';
  signal \-wp3\ : std_logic := '0';
  signal \-wp4\ : std_logic := '0';
  signal \-wp5\ : std_logic := '0';
  signal \-zero16.drive\ : std_logic := '0';
  signal \boot.trap\ : std_logic := '0';
  signal \bottom.1k\ : std_logic := '0';
  signal \bus.power.reset_l\ : std_logic := '0';
  signal \destimod0_l\ : std_logic := '0';
  signal \have_wrong_word\ : std_logic := '0';
  signal \inst_in_2nd_or_4th_quarter\ : std_logic := '0';
  signal \inst_in_left_half\ : std_logic := '0';
  signal \int.enable\ : std_logic := '0';
  signal \iwrited_l\ : std_logic := '0';
  signal \last_byte_in_word\ : std_logic := '0';
  signal \lc_byte_mode\ : std_logic := '0';
  signal \lm_drive_enb\ : std_logic := '0';
  signal \lpc.hold\ : std_logic := '0';
  signal \machruna_l\ : std_logic := '0';
  signal \mbusy.sync\ : std_logic := '0';
  signal \mempar_in\ : std_logic := '0';
  signal \mempar_out\ : std_logic := '0';
  signal \next.instr\ : std_logic := '0';
  signal \next.instrd\ : std_logic := '0';
  signal \pgf.or.int.or.sb\ : std_logic := '0';
  signal \pgf.or.int\ : std_logic := '0';
  signal \power_reset_a\ : std_logic := '0';
  signal \prog.boot\ : std_logic := '0';
  signal \prog.bus.reset\ : std_logic := '0';
  signal \prog.unibus.reset\ : std_logic := '0';
  signal \rd.in.progress\ : std_logic := '0';
  signal \sequence.break\ : std_logic := '0';
  signal \set.rd.in.progress\ : std_logic := '0';
  signal \stat.ovf\ : std_logic := '0';
  signal \use.md\ : std_logic := '0';
  signal \zero12.drive\ : std_logic := '0';
  signal \zero16.drive\ : std_logic := '0';
  signal a0 : std_logic := '0';
  signal a1 : std_logic := '0';
  signal a10 : std_logic := '0';
  signal a11 : std_logic := '0';
  signal a12 : std_logic := '0';
  signal a13 : std_logic := '0';
  signal a14 : std_logic := '0';
  signal a15 : std_logic := '0';
  signal a16 : std_logic := '0';
  signal a17 : std_logic := '0';
  signal a18 : std_logic := '0';
  signal a19 : std_logic := '0';
  signal a2 : std_logic := '0';
  signal a20 : std_logic := '0';
  signal a21 : std_logic := '0';
  signal a22 : std_logic := '0';
  signal a23 : std_logic := '0';
  signal a24 : std_logic := '0';
  signal a25 : std_logic := '0';
  signal a26 : std_logic := '0';
  signal a27 : std_logic := '0';
  signal a28 : std_logic := '0';
  signal a29 : std_logic := '0';
  signal a3 : std_logic := '0';
  signal a30 : std_logic := '0';
  signal a31a : std_logic := '0';
  signal a31b : std_logic := '0';
  signal a4 : std_logic := '0';
  signal a5 : std_logic := '0';
  signal a6 : std_logic := '0';
  signal a7 : std_logic := '0';
  signal a8 : std_logic := '0';
  signal a9 : std_logic := '0';
  signal aa0 : std_logic := '0';
  signal aa1 : std_logic := '0';
  signal aa10 : std_logic := '0';
  signal aa11 : std_logic := '0';
  signal aa12 : std_logic := '0';
  signal aa13 : std_logic := '0';
  signal aa14 : std_logic := '0';
  signal aa15 : std_logic := '0';
  signal aa16 : std_logic := '0';
  signal aa17 : std_logic := '0';
  signal aa2 : std_logic := '0';
  signal aa3 : std_logic := '0';
  signal aa4 : std_logic := '0';
  signal aa5 : std_logic := '0';
  signal aa6 : std_logic := '0';
  signal aa7 : std_logic := '0';
  signal aa8 : std_logic := '0';
  signal aa9 : std_logic := '0';
  signal aeqm : std_logic := '0';
  signal alu0 : std_logic := '0';
  signal alu1 : std_logic := '0';
  signal alu10 : std_logic := '0';
  signal alu11 : std_logic := '0';
  signal alu12 : std_logic := '0';
  signal alu13 : std_logic := '0';
  signal alu14 : std_logic := '0';
  signal alu15 : std_logic := '0';
  signal alu16 : std_logic := '0';
  signal alu17 : std_logic := '0';
  signal alu18 : std_logic := '0';
  signal alu19 : std_logic := '0';
  signal alu2 : std_logic := '0';
  signal alu20 : std_logic := '0';
  signal alu21 : std_logic := '0';
  signal alu22 : std_logic := '0';
  signal alu23 : std_logic := '0';
  signal alu24 : std_logic := '0';
  signal alu25 : std_logic := '0';
  signal alu26 : std_logic := '0';
  signal alu27 : std_logic := '0';
  signal alu28 : std_logic := '0';
  signal alu29 : std_logic := '0';
  signal alu3 : std_logic := '0';
  signal alu30 : std_logic := '0';
  signal alu31 : std_logic := '0';
  signal alu32 : std_logic := '0';
  signal alu4 : std_logic := '0';
  signal alu5 : std_logic := '0';
  signal alu6 : std_logic := '0';
  signal alu7 : std_logic := '0';
  signal alu8 : std_logic := '0';
  signal alu9 : std_logic := '0';
  signal aluadd : std_logic := '0';
  signal aluf0a : std_logic := '0';
  signal aluf0b : std_logic := '0';
  signal aluf1a : std_logic := '0';
  signal aluf1b : std_logic := '0';
  signal aluf2a : std_logic := '0';
  signal aluf2b : std_logic := '0';
  signal aluf3a : std_logic := '0';
  signal aluf3b : std_logic := '0';
  signal alumode : std_logic := '0';
  signal aluneg : std_logic := '0';
  signal alusub : std_logic := '0';
  signal amem0 : std_logic := '0';
  signal amem1 : std_logic := '0';
  signal amem10 : std_logic := '0';
  signal amem11 : std_logic := '0';
  signal amem12 : std_logic := '0';
  signal amem13 : std_logic := '0';
  signal amem14 : std_logic := '0';
  signal amem15 : std_logic := '0';
  signal amem16 : std_logic := '0';
  signal amem17 : std_logic := '0';
  signal amem18 : std_logic := '0';
  signal amem19 : std_logic := '0';
  signal amem2 : std_logic := '0';
  signal amem20 : std_logic := '0';
  signal amem21 : std_logic := '0';
  signal amem22 : std_logic := '0';
  signal amem23 : std_logic := '0';
  signal amem24 : std_logic := '0';
  signal amem25 : std_logic := '0';
  signal amem26 : std_logic := '0';
  signal amem27 : std_logic := '0';
  signal amem28 : std_logic := '0';
  signal amem29 : std_logic := '0';
  signal amem3 : std_logic := '0';
  signal amem30 : std_logic := '0';
  signal amem31 : std_logic := '0';
  signal amem4 : std_logic := '0';
  signal amem5 : std_logic := '0';
  signal amem6 : std_logic := '0';
  signal amem7 : std_logic := '0';
  signal amem8 : std_logic := '0';
  signal amem9 : std_logic := '0';
  signal amemparity : std_logic := '0';
  signal aparity : std_logic := '0';
  signal aparl : std_logic := '0';
  signal aparm : std_logic := '0';
  signal aparok : std_logic := '0';
  signal apass1 : std_logic := '0';
  signal apass2 : std_logic := '0';
  signal apassenb : std_logic := '0';
  signal clk1 : std_logic := '0';
  signal clk1a : std_logic := '0';
  signal clk2 : std_logic := '0';
  signal clk2a : std_logic := '0';
  signal clk2b : std_logic := '0';
  signal clk2c : std_logic := '0';
  signal clk3 : std_logic := '0';
  signal clk3a : std_logic := '0';
  signal clk3b : std_logic := '0';
  signal clk3c : std_logic := '0';
  signal clk3d : std_logic := '0';
  signal clk3e : std_logic := '0';
  signal clk3f : std_logic := '0';
  signal clk4 : std_logic := '0';
  signal clk4a : std_logic := '0';
  signal clk4b : std_logic := '0';
  signal clk4c : std_logic := '0';
  signal clk4d : std_logic := '0';
  signal clk4e : std_logic := '0';
  signal clk4f : std_logic := '0';
  signal clk5 : std_logic := '0';
  signal clk5a : std_logic := '0';
  signal conds0 : std_logic := '0';
  signal conds1 : std_logic := '0';
  signal conds2 : std_logic := '0';
  signal cyclecompleted : std_logic := '0';
  signal dadr10a : std_logic := '0';
  signal dadr10c : std_logic := '0';
  signal dc0 : std_logic := '0';
  signal dc1 : std_logic := '0';
  signal dc2 : std_logic := '0';
  signal dc3 : std_logic := '0';
  signal dc4 : std_logic := '0';
  signal dc5 : std_logic := '0';
  signal dc6 : std_logic := '0';
  signal dc7 : std_logic := '0';
  signal dc8 : std_logic := '0';
  signal dc9 : std_logic := '0';
  signal dcdrive : std_logic := '0';
  signal dest : std_logic := '0';
  signal destd : std_logic := '0';
  signal destm : std_logic := '0';
  signal destmd : std_logic := '0';
  signal destmdr : std_logic := '0';
  signal destmem : std_logic := '0';
  signal destspc : std_logic := '0';
  signal destspcd : std_logic := '0';
  signal dispenb : std_logic := '0';
  signal dispwr : std_logic := '0';
  signal divaddcond : std_logic := '0';
  signal divsubcond : std_logic := '0';
  signal dmask0 : std_logic := '0';
  signal dmask1 : std_logic := '0';
  signal dmask2 : std_logic := '0';
  signal dmask3 : std_logic := '0';
  signal dmask4 : std_logic := '0';
  signal dmask5 : std_logic := '0';
  signal dmask6 : std_logic := '0';
  signal dn : std_logic := '0';
  signal dp : std_logic := '0';
  signal dpar : std_logic := '0';
  signal dpareven : std_logic := '0';
  signal dparl : std_logic := '0';
  signal dparok : std_logic := '0';
  signal dpc0 : std_logic := '0';
  signal dpc1 : std_logic := '0';
  signal dpc10 : std_logic := '0';
  signal dpc11 : std_logic := '0';
  signal dpc12 : std_logic := '0';
  signal dpc13 : std_logic := '0';
  signal dpc2 : std_logic := '0';
  signal dpc3 : std_logic := '0';
  signal dpc4 : std_logic := '0';
  signal dpc5 : std_logic := '0';
  signal dpc6 : std_logic := '0';
  signal dpc7 : std_logic := '0';
  signal dpc8 : std_logic := '0';
  signal dpc9 : std_logic := '0';
  signal dpe : std_logic := '0';
  signal dr : std_logic := '0';
  signal eadr0 : std_logic := '0';
  signal eadr1 : std_logic := '0';
  signal eadr2 : std_logic := '0';
  signal eadr3 : std_logic := '0';
  signal err : std_logic := '0';
  signal errstop : std_logic := '0';
  signal gnd : std_logic := '0';
  signal hi1 : std_logic := '0';
  signal hi10 : std_logic := '0';
  signal hi11 : std_logic := '0';
  signal hi12 : std_logic := '0';
  signal hi2 : std_logic := '0';
  signal hi3 : std_logic := '0';
  signal hi4 : std_logic := '0';
  signal hi5 : std_logic := '0';
  signal hi6 : std_logic := '0';
  signal hi7 : std_logic := '0';
  signal hi8 : std_logic := '0';
  signal hi9 : std_logic := '0';
  signal highok : std_logic := '0';
  signal i0 : std_logic := '0';
  signal i1 : std_logic := '0';
  signal i10 : std_logic := '0';
  signal i11 : std_logic := '0';
  signal i12 : std_logic := '0';
  signal i13 : std_logic := '0';
  signal i14 : std_logic := '0';
  signal i15 : std_logic := '0';
  signal i16 : std_logic := '0';
  signal i17 : std_logic := '0';
  signal i18 : std_logic := '0';
  signal i19 : std_logic := '0';
  signal i2 : std_logic := '0';
  signal i20 : std_logic := '0';
  signal i21 : std_logic := '0';
  signal i22 : std_logic := '0';
  signal i23 : std_logic := '0';
  signal i24 : std_logic := '0';
  signal i25 : std_logic := '0';
  signal i26 : std_logic := '0';
  signal i27 : std_logic := '0';
  signal i28 : std_logic := '0';
  signal i29 : std_logic := '0';
  signal i3 : std_logic := '0';
  signal i30 : std_logic := '0';
  signal i31 : std_logic := '0';
  signal i32 : std_logic := '0';
  signal i33 : std_logic := '0';
  signal i34 : std_logic := '0';
  signal i35 : std_logic := '0';
  signal i36 : std_logic := '0';
  signal i37 : std_logic := '0';
  signal i38 : std_logic := '0';
  signal i39 : std_logic := '0';
  signal i4 : std_logic := '0';
  signal i40 : std_logic := '0';
  signal i41 : std_logic := '0';
  signal i42 : std_logic := '0';
  signal i43 : std_logic := '0';
  signal i44 : std_logic := '0';
  signal i45 : std_logic := '0';
  signal i46 : std_logic := '0';
  signal i47 : std_logic := '0';
  signal i48 : std_logic := '0';
  signal i5 : std_logic := '0';
  signal i6 : std_logic := '0';
  signal i7 : std_logic := '0';
  signal i8 : std_logic := '0';
  signal i9 : std_logic := '0';
  signal idebug : std_logic := '0';
  signal imod : std_logic := '0';
  signal imodd : std_logic := '0';
  signal inop : std_logic := '0';
  signal int : std_logic := '0';
  signal iob0 : std_logic := '0';
  signal iob1 : std_logic := '0';
  signal iob10 : std_logic := '0';
  signal iob11 : std_logic := '0';
  signal iob12 : std_logic := '0';
  signal iob13 : std_logic := '0';
  signal iob14 : std_logic := '0';
  signal iob15 : std_logic := '0';
  signal iob16 : std_logic := '0';
  signal iob17 : std_logic := '0';
  signal iob18 : std_logic := '0';
  signal iob19 : std_logic := '0';
  signal iob2 : std_logic := '0';
  signal iob20 : std_logic := '0';
  signal iob21 : std_logic := '0';
  signal iob22 : std_logic := '0';
  signal iob23 : std_logic := '0';
  signal iob24 : std_logic := '0';
  signal iob25 : std_logic := '0';
  signal iob26 : std_logic := '0';
  signal iob27 : std_logic := '0';
  signal iob28 : std_logic := '0';
  signal iob29 : std_logic := '0';
  signal iob3 : std_logic := '0';
  signal iob30 : std_logic := '0';
  signal iob31 : std_logic := '0';
  signal iob32 : std_logic := '0';
  signal iob33 : std_logic := '0';
  signal iob34 : std_logic := '0';
  signal iob35 : std_logic := '0';
  signal iob36 : std_logic := '0';
  signal iob37 : std_logic := '0';
  signal iob38 : std_logic := '0';
  signal iob39 : std_logic := '0';
  signal iob4 : std_logic := '0';
  signal iob40 : std_logic := '0';
  signal iob41 : std_logic := '0';
  signal iob42 : std_logic := '0';
  signal iob43 : std_logic := '0';
  signal iob44 : std_logic := '0';
  signal iob45 : std_logic := '0';
  signal iob46 : std_logic := '0';
  signal iob47 : std_logic := '0';
  signal iob5 : std_logic := '0';
  signal iob6 : std_logic := '0';
  signal iob7 : std_logic := '0';
  signal iob8 : std_logic := '0';
  signal iob9 : std_logic := '0';
  signal ipar0 : std_logic := '0';
  signal ipar1 : std_logic := '0';
  signal ipar2 : std_logic := '0';
  signal ipar3 : std_logic := '0';
  signal iparity : std_logic := '0';
  signal iparok : std_logic := '0';
  signal ipc0 : std_logic := '0';
  signal ipc1 : std_logic := '0';
  signal ipc10 : std_logic := '0';
  signal ipc11 : std_logic := '0';
  signal ipc12 : std_logic := '0';
  signal ipc13 : std_logic := '0';
  signal ipc2 : std_logic := '0';
  signal ipc3 : std_logic := '0';
  signal ipc4 : std_logic := '0';
  signal ipc5 : std_logic := '0';
  signal ipc6 : std_logic := '0';
  signal ipc7 : std_logic := '0';
  signal ipc8 : std_logic := '0';
  signal ipc9 : std_logic := '0';
  signal ipe : std_logic := '0';
  signal ir0 : std_logic := '0';
  signal ir1 : std_logic := '0';
  signal ir10 : std_logic := '0';
  signal ir11 : std_logic := '0';
  signal ir12 : std_logic := '0';
  signal ir12b : std_logic := '0';
  signal ir13 : std_logic := '0';
  signal ir13b : std_logic := '0';
  signal ir14 : std_logic := '0';
  signal ir14b : std_logic := '0';
  signal ir15 : std_logic := '0';
  signal ir15b : std_logic := '0';
  signal ir16 : std_logic := '0';
  signal ir16b : std_logic := '0';
  signal ir17 : std_logic := '0';
  signal ir17b : std_logic := '0';
  signal ir18 : std_logic := '0';
  signal ir18b : std_logic := '0';
  signal ir19 : std_logic := '0';
  signal ir19b : std_logic := '0';
  signal ir2 : std_logic := '0';
  signal ir20 : std_logic := '0';
  signal ir20b : std_logic := '0';
  signal ir21 : std_logic := '0';
  signal ir21b : std_logic := '0';
  signal ir22 : std_logic := '0';
  signal ir22b : std_logic := '0';
  signal ir23 : std_logic := '0';
  signal ir24 : std_logic := '0';
  signal ir25 : std_logic := '0';
  signal ir26 : std_logic := '0';
  signal ir27 : std_logic := '0';
  signal ir28 : std_logic := '0';
  signal ir29 : std_logic := '0';
  signal ir3 : std_logic := '0';
  signal ir30 : std_logic := '0';
  signal ir31 : std_logic := '0';
  signal ir32 : std_logic := '0';
  signal ir33 : std_logic := '0';
  signal ir34 : std_logic := '0';
  signal ir35 : std_logic := '0';
  signal ir36 : std_logic := '0';
  signal ir37 : std_logic := '0';
  signal ir38 : std_logic := '0';
  signal ir39 : std_logic := '0';
  signal ir4 : std_logic := '0';
  signal ir40 : std_logic := '0';
  signal ir41 : std_logic := '0';
  signal ir42 : std_logic := '0';
  signal ir43 : std_logic := '0';
  signal ir44 : std_logic := '0';
  signal ir45 : std_logic := '0';
  signal ir46 : std_logic := '0';
  signal ir47 : std_logic := '0';
  signal ir48 : std_logic := '0';
  signal ir5 : std_logic := '0';
  signal ir6 : std_logic := '0';
  signal ir7 : std_logic := '0';
  signal ir8 : std_logic := '0';
  signal ir8b : std_logic := '0';
  signal ir9 : std_logic := '0';
  signal ir9b : std_logic := '0';
  signal iralu : std_logic := '0';
  signal irdisp : std_logic := '0';
  signal irjump : std_logic := '0';
  signal iwr0 : std_logic := '0';
  signal iwr1 : std_logic := '0';
  signal iwr10 : std_logic := '0';
  signal iwr11 : std_logic := '0';
  signal iwr12 : std_logic := '0';
  signal iwr13 : std_logic := '0';
  signal iwr14 : std_logic := '0';
  signal iwr15 : std_logic := '0';
  signal iwr16 : std_logic := '0';
  signal iwr17 : std_logic := '0';
  signal iwr18 : std_logic := '0';
  signal iwr19 : std_logic := '0';
  signal iwr2 : std_logic := '0';
  signal iwr20 : std_logic := '0';
  signal iwr21 : std_logic := '0';
  signal iwr22 : std_logic := '0';
  signal iwr23 : std_logic := '0';
  signal iwr24 : std_logic := '0';
  signal iwr25 : std_logic := '0';
  signal iwr26 : std_logic := '0';
  signal iwr27 : std_logic := '0';
  signal iwr28 : std_logic := '0';
  signal iwr29 : std_logic := '0';
  signal iwr3 : std_logic := '0';
  signal iwr30 : std_logic := '0';
  signal iwr31 : std_logic := '0';
  signal iwr32 : std_logic := '0';
  signal iwr33 : std_logic := '0';
  signal iwr34 : std_logic := '0';
  signal iwr35 : std_logic := '0';
  signal iwr36 : std_logic := '0';
  signal iwr37 : std_logic := '0';
  signal iwr38 : std_logic := '0';
  signal iwr39 : std_logic := '0';
  signal iwr4 : std_logic := '0';
  signal iwr40 : std_logic := '0';
  signal iwr41 : std_logic := '0';
  signal iwr42 : std_logic := '0';
  signal iwr43 : std_logic := '0';
  signal iwr44 : std_logic := '0';
  signal iwr45 : std_logic := '0';
  signal iwr46 : std_logic := '0';
  signal iwr47 : std_logic := '0';
  signal iwr48 : std_logic := '0';
  signal iwr5 : std_logic := '0';
  signal iwr6 : std_logic := '0';
  signal iwr7 : std_logic := '0';
  signal iwr8 : std_logic := '0';
  signal iwr9 : std_logic := '0';
  signal iwrite : std_logic := '0';
  signal iwrited : std_logic := '0';
  signal iwriteda : std_logic := '0';
  signal iwritedb : std_logic := '0';
  signal iwritedc : std_logic := '0';
  signal iwritedd : std_logic := '0';
  signal iwrp1 : std_logic := '0';
  signal iwrp2 : std_logic := '0';
  signal iwrp3 : std_logic := '0';
  signal iwrp4 : std_logic := '0';
  signal jcalf : std_logic := '0';
  signal jcond : std_logic := '0';
  signal jfalse : std_logic := '0';
  signal jret : std_logic := '0';
  signal jretf : std_logic := '0';
  signal l0 : std_logic := '0';
  signal l1 : std_logic := '0';
  signal l10 : std_logic := '0';
  signal l11 : std_logic := '0';
  signal l12 : std_logic := '0';
  signal l13 : std_logic := '0';
  signal l14 : std_logic := '0';
  signal l15 : std_logic := '0';
  signal l16 : std_logic := '0';
  signal l17 : std_logic := '0';
  signal l18 : std_logic := '0';
  signal l19 : std_logic := '0';
  signal l2 : std_logic := '0';
  signal l20 : std_logic := '0';
  signal l21 : std_logic := '0';
  signal l22 : std_logic := '0';
  signal l23 : std_logic := '0';
  signal l24 : std_logic := '0';
  signal l25 : std_logic := '0';
  signal l26 : std_logic := '0';
  signal l27 : std_logic := '0';
  signal l28 : std_logic := '0';
  signal l29 : std_logic := '0';
  signal l3 : std_logic := '0';
  signal l30 : std_logic := '0';
  signal l31 : std_logic := '0';
  signal l4 : std_logic := '0';
  signal l5 : std_logic := '0';
  signal l6 : std_logic := '0';
  signal l7 : std_logic := '0';
  signal l8 : std_logic := '0';
  signal l9 : std_logic := '0';
  signal lc0 : std_logic := '0';
  signal lc0b : std_logic := '0';
  signal lc1 : std_logic := '0';
  signal lc10 : std_logic := '0';
  signal lc11 : std_logic := '0';
  signal lc12 : std_logic := '0';
  signal lc13 : std_logic := '0';
  signal lc14 : std_logic := '0';
  signal lc15 : std_logic := '0';
  signal lc16 : std_logic := '0';
  signal lc17 : std_logic := '0';
  signal lc18 : std_logic := '0';
  signal lc19 : std_logic := '0';
  signal lc2 : std_logic := '0';
  signal lc20 : std_logic := '0';
  signal lc21 : std_logic := '0';
  signal lc22 : std_logic := '0';
  signal lc23 : std_logic := '0';
  signal lc24 : std_logic := '0';
  signal lc25 : std_logic := '0';
  signal lc3 : std_logic := '0';
  signal lc4 : std_logic := '0';
  signal lc5 : std_logic := '0';
  signal lc6 : std_logic := '0';
  signal lc7 : std_logic := '0';
  signal lc8 : std_logic := '0';
  signal lc9 : std_logic := '0';
  signal lca0 : std_logic := '0';
  signal lca1 : std_logic := '0';
  signal lca2 : std_logic := '0';
  signal lca3 : std_logic := '0';
  signal lcdrive : std_logic := '0';
  signal lcinc : std_logic := '0';
  signal lcry3 : std_logic := '0';
  signal ldmode : std_logic := '0';
  signal ldstat : std_logic := '0';
  signal loadmd : std_logic := '0';
  signal lparity : std_logic := '0';
  signal lparl : std_logic := '0';
  signal lpc0 : std_logic := '0';
  signal lpc1 : std_logic := '0';
  signal lpc10 : std_logic := '0';
  signal lpc11 : std_logic := '0';
  signal lpc12 : std_logic := '0';
  signal lpc13 : std_logic := '0';
  signal lpc2 : std_logic := '0';
  signal lpc3 : std_logic := '0';
  signal lpc4 : std_logic := '0';
  signal lpc5 : std_logic := '0';
  signal lpc6 : std_logic := '0';
  signal lpc7 : std_logic := '0';
  signal lpc8 : std_logic := '0';
  signal lpc9 : std_logic := '0';
  signal m0 : std_logic := '0';
  signal m1 : std_logic := '0';
  signal m10 : std_logic := '0';
  signal m11 : std_logic := '0';
  signal m12 : std_logic := '0';
  signal m13 : std_logic := '0';
  signal m14 : std_logic := '0';
  signal m15 : std_logic := '0';
  signal m16 : std_logic := '0';
  signal m17 : std_logic := '0';
  signal m18 : std_logic := '0';
  signal m19 : std_logic := '0';
  signal m2 : std_logic := '0';
  signal m20 : std_logic := '0';
  signal m21 : std_logic := '0';
  signal m22 : std_logic := '0';
  signal m23 : std_logic := '0';
  signal m24 : std_logic := '0';
  signal m25 : std_logic := '0';
  signal m26 : std_logic := '0';
  signal m27 : std_logic := '0';
  signal m28 : std_logic := '0';
  signal m29 : std_logic := '0';
  signal m3 : std_logic := '0';
  signal m30 : std_logic := '0';
  signal m31 : std_logic := '0';
  signal m31b : std_logic := '0';
  signal m4 : std_logic := '0';
  signal m5 : std_logic := '0';
  signal m6 : std_logic := '0';
  signal m7 : std_logic := '0';
  signal m8 : std_logic := '0';
  signal m9 : std_logic := '0';
  signal machrun : std_logic := '0';
  signal mapi10 : std_logic := '0';
  signal mapi11 : std_logic := '0';
  signal mapi12 : std_logic := '0';
  signal mapi13 : std_logic := '0';
  signal mapi14 : std_logic := '0';
  signal mapi15 : std_logic := '0';
  signal mapi16 : std_logic := '0';
  signal mapi17 : std_logic := '0';
  signal mapi18 : std_logic := '0';
  signal mapi19 : std_logic := '0';
  signal mapi20 : std_logic := '0';
  signal mapi21 : std_logic := '0';
  signal mapi22 : std_logic := '0';
  signal mapi23 : std_logic := '0';
  signal mapi8 : std_logic := '0';
  signal mapi9 : std_logic := '0';
  signal mapwr0d : std_logic := '0';
  signal mapwr1d : std_logic := '0';
  signal mbusy : std_logic := '0';
  signal mclk1 : std_logic := '0';
  signal mclk1a : std_logic := '0';
  signal mclk5 : std_logic := '0';
  signal mclk5a : std_logic := '0';
  signal mclk7 : std_logic := '0';
  signal mdclk : std_logic := '0';
  signal mdgetspar : std_logic := '0';
  signal mdhaspar : std_logic := '0';
  signal mdpar : std_logic := '0';
  signal mdparerr : std_logic := '0';
  signal mdpareven : std_logic := '0';
  signal mdparl : std_logic := '0';
  signal mdparm : std_logic := '0';
  signal mdparodd : std_logic := '0';
  signal mdsela : std_logic := '0';
  signal mdselb : std_logic := '0';
  signal mem0 : std_logic := '0';
  signal mem1 : std_logic := '0';
  signal mem10 : std_logic := '0';
  signal mem11 : std_logic := '0';
  signal mem12 : std_logic := '0';
  signal mem13 : std_logic := '0';
  signal mem14 : std_logic := '0';
  signal mem15 : std_logic := '0';
  signal mem16 : std_logic := '0';
  signal mem17 : std_logic := '0';
  signal mem18 : std_logic := '0';
  signal mem19 : std_logic := '0';
  signal mem2 : std_logic := '0';
  signal mem20 : std_logic := '0';
  signal mem21 : std_logic := '0';
  signal mem22 : std_logic := '0';
  signal mem23 : std_logic := '0';
  signal mem24 : std_logic := '0';
  signal mem25 : std_logic := '0';
  signal mem26 : std_logic := '0';
  signal mem27 : std_logic := '0';
  signal mem28 : std_logic := '0';
  signal mem29 : std_logic := '0';
  signal mem3 : std_logic := '0';
  signal mem30 : std_logic := '0';
  signal mem31 : std_logic := '0';
  signal mem4 : std_logic := '0';
  signal mem5 : std_logic := '0';
  signal mem6 : std_logic := '0';
  signal mem7 : std_logic := '0';
  signal mem8 : std_logic := '0';
  signal mem9 : std_logic := '0';
  signal memparok : std_logic := '0';
  signal memprepare : std_logic := '0';
  signal memrq : std_logic := '0';
  signal memstart : std_logic := '0';
  signal mf0 : std_logic := '0';
  signal mf1 : std_logic := '0';
  signal mf10 : std_logic := '0';
  signal mf11 : std_logic := '0';
  signal mf12 : std_logic := '0';
  signal mf13 : std_logic := '0';
  signal mf14 : std_logic := '0';
  signal mf15 : std_logic := '0';
  signal mf16 : std_logic := '0';
  signal mf17 : std_logic := '0';
  signal mf18 : std_logic := '0';
  signal mf19 : std_logic := '0';
  signal mf2 : std_logic := '0';
  signal mf20 : std_logic := '0';
  signal mf21 : std_logic := '0';
  signal mf22 : std_logic := '0';
  signal mf23 : std_logic := '0';
  signal mf24 : std_logic := '0';
  signal mf25 : std_logic := '0';
  signal mf26 : std_logic := '0';
  signal mf27 : std_logic := '0';
  signal mf28 : std_logic := '0';
  signal mf29 : std_logic := '0';
  signal mf3 : std_logic := '0';
  signal mf30 : std_logic := '0';
  signal mf31 : std_logic := '0';
  signal mf4 : std_logic := '0';
  signal mf5 : std_logic := '0';
  signal mf6 : std_logic := '0';
  signal mf7 : std_logic := '0';
  signal mf8 : std_logic := '0';
  signal mf9 : std_logic := '0';
  signal mfdrive : std_logic := '0';
  signal mfenb : std_logic := '0';
  signal mmem0 : std_logic := '0';
  signal mmem1 : std_logic := '0';
  signal mmem10 : std_logic := '0';
  signal mmem11 : std_logic := '0';
  signal mmem12 : std_logic := '0';
  signal mmem13 : std_logic := '0';
  signal mmem14 : std_logic := '0';
  signal mmem15 : std_logic := '0';
  signal mmem16 : std_logic := '0';
  signal mmem17 : std_logic := '0';
  signal mmem18 : std_logic := '0';
  signal mmem19 : std_logic := '0';
  signal mmem2 : std_logic := '0';
  signal mmem20 : std_logic := '0';
  signal mmem21 : std_logic := '0';
  signal mmem22 : std_logic := '0';
  signal mmem23 : std_logic := '0';
  signal mmem24 : std_logic := '0';
  signal mmem25 : std_logic := '0';
  signal mmem26 : std_logic := '0';
  signal mmem27 : std_logic := '0';
  signal mmem28 : std_logic := '0';
  signal mmem29 : std_logic := '0';
  signal mmem3 : std_logic := '0';
  signal mmem30 : std_logic := '0';
  signal mmem31 : std_logic := '0';
  signal mmem4 : std_logic := '0';
  signal mmem5 : std_logic := '0';
  signal mmem6 : std_logic := '0';
  signal mmem7 : std_logic := '0';
  signal mmem8 : std_logic := '0';
  signal mmem9 : std_logic := '0';
  signal mmemparity : std_logic := '0';
  signal mmemparok : std_logic := '0';
  signal mpareven : std_logic := '0';
  signal mparity : std_logic := '0';
  signal mparl : std_logic := '0';
  signal mparm : std_logic := '0';
  signal mparodd : std_logic := '0';
  signal mpass : std_logic := '0';
  signal mpassl : std_logic := '0';
  signal msk0 : std_logic := '0';
  signal msk1 : std_logic := '0';
  signal msk10 : std_logic := '0';
  signal msk11 : std_logic := '0';
  signal msk12 : std_logic := '0';
  signal msk13 : std_logic := '0';
  signal msk14 : std_logic := '0';
  signal msk15 : std_logic := '0';
  signal msk16 : std_logic := '0';
  signal msk17 : std_logic := '0';
  signal msk18 : std_logic := '0';
  signal msk19 : std_logic := '0';
  signal msk2 : std_logic := '0';
  signal msk20 : std_logic := '0';
  signal msk21 : std_logic := '0';
  signal msk22 : std_logic := '0';
  signal msk23 : std_logic := '0';
  signal msk24 : std_logic := '0';
  signal msk25 : std_logic := '0';
  signal msk26 : std_logic := '0';
  signal msk27 : std_logic := '0';
  signal msk28 : std_logic := '0';
  signal msk29 : std_logic := '0';
  signal msk3 : std_logic := '0';
  signal msk30 : std_logic := '0';
  signal msk31 : std_logic := '0';
  signal msk4 : std_logic := '0';
  signal msk5 : std_logic := '0';
  signal msk6 : std_logic := '0';
  signal msk7 : std_logic := '0';
  signal msk8 : std_logic := '0';
  signal msk9 : std_logic := '0';
  signal mskl0 : std_logic := '0';
  signal mskl1 : std_logic := '0';
  signal mskl2 : std_logic := '0';
  signal mskl3 : std_logic := '0';
  signal mskl3cry : std_logic := '0';
  signal mskl4 : std_logic := '0';
  signal mskr0 : std_logic := '0';
  signal mskr1 : std_logic := '0';
  signal mskr2 : std_logic := '0';
  signal mskr3 : std_logic := '0';
  signal mskr4 : std_logic := '0';
  signal n : std_logic := '0';
  signal needfetch : std_logic := '0';
  signal newlc : std_logic := '0';
  signal nop : std_logic := '0';
  signal nop11 : std_logic := '0';
  signal nopa : std_logic := '0';
  signal npc0 : std_logic := '0';
  signal npc1 : std_logic := '0';
  signal npc10 : std_logic := '0';
  signal npc11 : std_logic := '0';
  signal npc12 : std_logic := '0';
  signal npc13 : std_logic := '0';
  signal npc2 : std_logic := '0';
  signal npc3 : std_logic := '0';
  signal npc4 : std_logic := '0';
  signal npc5 : std_logic := '0';
  signal npc6 : std_logic := '0';
  signal npc7 : std_logic := '0';
  signal npc8 : std_logic := '0';
  signal npc9 : std_logic := '0';
  signal ob0 : std_logic := '0';
  signal ob1 : std_logic := '0';
  signal ob10 : std_logic := '0';
  signal ob11 : std_logic := '0';
  signal ob12 : std_logic := '0';
  signal ob13 : std_logic := '0';
  signal ob14 : std_logic := '0';
  signal ob15 : std_logic := '0';
  signal ob16 : std_logic := '0';
  signal ob17 : std_logic := '0';
  signal ob18 : std_logic := '0';
  signal ob19 : std_logic := '0';
  signal ob2 : std_logic := '0';
  signal ob20 : std_logic := '0';
  signal ob21 : std_logic := '0';
  signal ob22 : std_logic := '0';
  signal ob23 : std_logic := '0';
  signal ob24 : std_logic := '0';
  signal ob25 : std_logic := '0';
  signal ob26 : std_logic := '0';
  signal ob27 : std_logic := '0';
  signal ob28 : std_logic := '0';
  signal ob29 : std_logic := '0';
  signal ob3 : std_logic := '0';
  signal ob30 : std_logic := '0';
  signal ob31 : std_logic := '0';
  signal ob4 : std_logic := '0';
  signal ob5 : std_logic := '0';
  signal ob6 : std_logic := '0';
  signal ob7 : std_logic := '0';
  signal ob8 : std_logic := '0';
  signal ob9 : std_logic := '0';
  signal opc0 : std_logic := '0';
  signal opc1 : std_logic := '0';
  signal opc10 : std_logic := '0';
  signal opc11 : std_logic := '0';
  signal opc12 : std_logic := '0';
  signal opc13 : std_logic := '0';
  signal opc2 : std_logic := '0';
  signal opc3 : std_logic := '0';
  signal opc4 : std_logic := '0';
  signal opc5 : std_logic := '0';
  signal opc6 : std_logic := '0';
  signal opc7 : std_logic := '0';
  signal opc8 : std_logic := '0';
  signal opc9 : std_logic := '0';
  signal opcclk : std_logic := '0';
  signal opcclka : std_logic := '0';
  signal opcclkb : std_logic := '0';
  signal opcclkc : std_logic := '0';
  signal opcinh : std_logic := '0';
  signal opcinha : std_logic := '0';
  signal opcinhb : std_logic := '0';
  signal osel0a : std_logic := '0';
  signal osel0b : std_logic := '0';
  signal osel1a : std_logic := '0';
  signal osel1b : std_logic := '0';
  signal pc0 : std_logic := '0';
  signal pc0a : std_logic := '0';
  signal pc0b : std_logic := '0';
  signal pc0c : std_logic := '0';
  signal pc0d : std_logic := '0';
  signal pc0e : std_logic := '0';
  signal pc0f : std_logic := '0';
  signal pc0g : std_logic := '0';
  signal pc0h : std_logic := '0';
  signal pc0i : std_logic := '0';
  signal pc0j : std_logic := '0';
  signal pc0k : std_logic := '0';
  signal pc0l : std_logic := '0';
  signal pc0m : std_logic := '0';
  signal pc0n : std_logic := '0';
  signal pc0o : std_logic := '0';
  signal pc0p : std_logic := '0';
  signal pc1 : std_logic := '0';
  signal pc10 : std_logic := '0';
  signal pc10a : std_logic := '0';
  signal pc10b : std_logic := '0';
  signal pc10c : std_logic := '0';
  signal pc10d : std_logic := '0';
  signal pc10e : std_logic := '0';
  signal pc10f : std_logic := '0';
  signal pc10g : std_logic := '0';
  signal pc10h : std_logic := '0';
  signal pc10i : std_logic := '0';
  signal pc10j : std_logic := '0';
  signal pc10k : std_logic := '0';
  signal pc10l : std_logic := '0';
  signal pc10m : std_logic := '0';
  signal pc10n : std_logic := '0';
  signal pc10o : std_logic := '0';
  signal pc10p : std_logic := '0';
  signal pc11 : std_logic := '0';
  signal pc11a : std_logic := '0';
  signal pc11b : std_logic := '0';
  signal pc11c : std_logic := '0';
  signal pc11d : std_logic := '0';
  signal pc11e : std_logic := '0';
  signal pc11f : std_logic := '0';
  signal pc11g : std_logic := '0';
  signal pc11h : std_logic := '0';
  signal pc11i : std_logic := '0';
  signal pc11j : std_logic := '0';
  signal pc11k : std_logic := '0';
  signal pc11l : std_logic := '0';
  signal pc11m : std_logic := '0';
  signal pc11n : std_logic := '0';
  signal pc11o : std_logic := '0';
  signal pc11p : std_logic := '0';
  signal pc12 : std_logic := '0';
  signal pc12b : std_logic := '0';
  signal pc13 : std_logic := '0';
  signal pc13b : std_logic := '0';
  signal pc1a : std_logic := '0';
  signal pc1b : std_logic := '0';
  signal pc1c : std_logic := '0';
  signal pc1d : std_logic := '0';
  signal pc1e : std_logic := '0';
  signal pc1f : std_logic := '0';
  signal pc1g : std_logic := '0';
  signal pc1h : std_logic := '0';
  signal pc1i : std_logic := '0';
  signal pc1j : std_logic := '0';
  signal pc1k : std_logic := '0';
  signal pc1l : std_logic := '0';
  signal pc1m : std_logic := '0';
  signal pc1n : std_logic := '0';
  signal pc1o : std_logic := '0';
  signal pc1p : std_logic := '0';
  signal pc2 : std_logic := '0';
  signal pc2a : std_logic := '0';
  signal pc2b : std_logic := '0';
  signal pc2c : std_logic := '0';
  signal pc2d : std_logic := '0';
  signal pc2e : std_logic := '0';
  signal pc2f : std_logic := '0';
  signal pc2g : std_logic := '0';
  signal pc2h : std_logic := '0';
  signal pc2i : std_logic := '0';
  signal pc2j : std_logic := '0';
  signal pc2k : std_logic := '0';
  signal pc2l : std_logic := '0';
  signal pc2m : std_logic := '0';
  signal pc2n : std_logic := '0';
  signal pc2o : std_logic := '0';
  signal pc2p : std_logic := '0';
  signal pc3 : std_logic := '0';
  signal pc3a : std_logic := '0';
  signal pc3b : std_logic := '0';
  signal pc3c : std_logic := '0';
  signal pc3d : std_logic := '0';
  signal pc3e : std_logic := '0';
  signal pc3f : std_logic := '0';
  signal pc3g : std_logic := '0';
  signal pc3h : std_logic := '0';
  signal pc3i : std_logic := '0';
  signal pc3j : std_logic := '0';
  signal pc3k : std_logic := '0';
  signal pc3l : std_logic := '0';
  signal pc3m : std_logic := '0';
  signal pc3n : std_logic := '0';
  signal pc3o : std_logic := '0';
  signal pc3p : std_logic := '0';
  signal pc4 : std_logic := '0';
  signal pc4a : std_logic := '0';
  signal pc4b : std_logic := '0';
  signal pc4c : std_logic := '0';
  signal pc4d : std_logic := '0';
  signal pc4e : std_logic := '0';
  signal pc4f : std_logic := '0';
  signal pc4g : std_logic := '0';
  signal pc4h : std_logic := '0';
  signal pc4i : std_logic := '0';
  signal pc4j : std_logic := '0';
  signal pc4k : std_logic := '0';
  signal pc4l : std_logic := '0';
  signal pc4m : std_logic := '0';
  signal pc4n : std_logic := '0';
  signal pc4o : std_logic := '0';
  signal pc4p : std_logic := '0';
  signal pc5 : std_logic := '0';
  signal pc5a : std_logic := '0';
  signal pc5b : std_logic := '0';
  signal pc5c : std_logic := '0';
  signal pc5d : std_logic := '0';
  signal pc5e : std_logic := '0';
  signal pc5f : std_logic := '0';
  signal pc5g : std_logic := '0';
  signal pc5h : std_logic := '0';
  signal pc5i : std_logic := '0';
  signal pc5j : std_logic := '0';
  signal pc5k : std_logic := '0';
  signal pc5l : std_logic := '0';
  signal pc5m : std_logic := '0';
  signal pc5n : std_logic := '0';
  signal pc5o : std_logic := '0';
  signal pc5p : std_logic := '0';
  signal pc6 : std_logic := '0';
  signal pc6a : std_logic := '0';
  signal pc6b : std_logic := '0';
  signal pc6c : std_logic := '0';
  signal pc6d : std_logic := '0';
  signal pc6e : std_logic := '0';
  signal pc6f : std_logic := '0';
  signal pc6g : std_logic := '0';
  signal pc6h : std_logic := '0';
  signal pc6i : std_logic := '0';
  signal pc6j : std_logic := '0';
  signal pc6k : std_logic := '0';
  signal pc6l : std_logic := '0';
  signal pc6m : std_logic := '0';
  signal pc6n : std_logic := '0';
  signal pc6o : std_logic := '0';
  signal pc6p : std_logic := '0';
  signal pc7 : std_logic := '0';
  signal pc7a : std_logic := '0';
  signal pc7b : std_logic := '0';
  signal pc7c : std_logic := '0';
  signal pc7d : std_logic := '0';
  signal pc7e : std_logic := '0';
  signal pc7f : std_logic := '0';
  signal pc7g : std_logic := '0';
  signal pc7h : std_logic := '0';
  signal pc7i : std_logic := '0';
  signal pc7j : std_logic := '0';
  signal pc7k : std_logic := '0';
  signal pc7l : std_logic := '0';
  signal pc7m : std_logic := '0';
  signal pc7n : std_logic := '0';
  signal pc7o : std_logic := '0';
  signal pc7p : std_logic := '0';
  signal pc8 : std_logic := '0';
  signal pc8a : std_logic := '0';
  signal pc8b : std_logic := '0';
  signal pc8c : std_logic := '0';
  signal pc8d : std_logic := '0';
  signal pc8e : std_logic := '0';
  signal pc8f : std_logic := '0';
  signal pc8g : std_logic := '0';
  signal pc8h : std_logic := '0';
  signal pc8i : std_logic := '0';
  signal pc8j : std_logic := '0';
  signal pc8k : std_logic := '0';
  signal pc8l : std_logic := '0';
  signal pc8m : std_logic := '0';
  signal pc8n : std_logic := '0';
  signal pc8o : std_logic := '0';
  signal pc8p : std_logic := '0';
  signal pc9 : std_logic := '0';
  signal pc9a : std_logic := '0';
  signal pc9b : std_logic := '0';
  signal pc9c : std_logic := '0';
  signal pc9d : std_logic := '0';
  signal pc9e : std_logic := '0';
  signal pc9f : std_logic := '0';
  signal pc9g : std_logic := '0';
  signal pc9h : std_logic := '0';
  signal pc9i : std_logic := '0';
  signal pc9j : std_logic := '0';
  signal pc9k : std_logic := '0';
  signal pc9l : std_logic := '0';
  signal pc9m : std_logic := '0';
  signal pc9n : std_logic := '0';
  signal pc9o : std_logic := '0';
  signal pc9p : std_logic := '0';
  signal pccry11 : std_logic := '0';
  signal pccry3 : std_logic := '0';
  signal pccry7 : std_logic := '0';
  signal pcs0 : std_logic := '0';
  signal pcs1 : std_logic := '0';
  signal pdl0 : std_logic := '0';
  signal pdl1 : std_logic := '0';
  signal pdl10 : std_logic := '0';
  signal pdl11 : std_logic := '0';
  signal pdl12 : std_logic := '0';
  signal pdl13 : std_logic := '0';
  signal pdl14 : std_logic := '0';
  signal pdl15 : std_logic := '0';
  signal pdl16 : std_logic := '0';
  signal pdl17 : std_logic := '0';
  signal pdl18 : std_logic := '0';
  signal pdl19 : std_logic := '0';
  signal pdl2 : std_logic := '0';
  signal pdl20 : std_logic := '0';
  signal pdl21 : std_logic := '0';
  signal pdl22 : std_logic := '0';
  signal pdl23 : std_logic := '0';
  signal pdl24 : std_logic := '0';
  signal pdl25 : std_logic := '0';
  signal pdl26 : std_logic := '0';
  signal pdl27 : std_logic := '0';
  signal pdl28 : std_logic := '0';
  signal pdl29 : std_logic := '0';
  signal pdl3 : std_logic := '0';
  signal pdl30 : std_logic := '0';
  signal pdl31 : std_logic := '0';
  signal pdl4 : std_logic := '0';
  signal pdl5 : std_logic := '0';
  signal pdl6 : std_logic := '0';
  signal pdl7 : std_logic := '0';
  signal pdl8 : std_logic := '0';
  signal pdl9 : std_logic := '0';
  signal pdlenb : std_logic := '0';
  signal pdlidx0 : std_logic := '0';
  signal pdlidx1 : std_logic := '0';
  signal pdlidx2 : std_logic := '0';
  signal pdlidx3 : std_logic := '0';
  signal pdlidx4 : std_logic := '0';
  signal pdlidx5 : std_logic := '0';
  signal pdlidx6 : std_logic := '0';
  signal pdlidx7 : std_logic := '0';
  signal pdlidx8 : std_logic := '0';
  signal pdlidx9 : std_logic := '0';
  signal pdlparity : std_logic := '0';
  signal pdlparok : std_logic := '0';
  signal pdlptr0 : std_logic := '0';
  signal pdlptr1 : std_logic := '0';
  signal pdlptr2 : std_logic := '0';
  signal pdlptr3 : std_logic := '0';
  signal pdlptr4 : std_logic := '0';
  signal pdlptr5 : std_logic := '0';
  signal pdlptr6 : std_logic := '0';
  signal pdlptr7 : std_logic := '0';
  signal pdlptr8 : std_logic := '0';
  signal pdlptr9 : std_logic := '0';
  signal pdlwrite : std_logic := '0';
  signal pdlwrited : std_logic := '0';
  signal pidrive : std_logic := '0';
  signal popj : std_logic := '0';
  signal promdisable : std_logic := '0';
  signal promdisabled : std_logic := '0';
  signal promenable : std_logic := '0';
  signal pwidx : std_logic := '0';
  signal q0 : std_logic := '0';
  signal q1 : std_logic := '0';
  signal q10 : std_logic := '0';
  signal q11 : std_logic := '0';
  signal q12 : std_logic := '0';
  signal q13 : std_logic := '0';
  signal q14 : std_logic := '0';
  signal q15 : std_logic := '0';
  signal q16 : std_logic := '0';
  signal q17 : std_logic := '0';
  signal q18 : std_logic := '0';
  signal q19 : std_logic := '0';
  signal q2 : std_logic := '0';
  signal q20 : std_logic := '0';
  signal q21 : std_logic := '0';
  signal q22 : std_logic := '0';
  signal q23 : std_logic := '0';
  signal q24 : std_logic := '0';
  signal q25 : std_logic := '0';
  signal q26 : std_logic := '0';
  signal q27 : std_logic := '0';
  signal q28 : std_logic := '0';
  signal q29 : std_logic := '0';
  signal q3 : std_logic := '0';
  signal q30 : std_logic := '0';
  signal q31 : std_logic := '0';
  signal q4 : std_logic := '0';
  signal q5 : std_logic := '0';
  signal q6 : std_logic := '0';
  signal q7 : std_logic := '0';
  signal q8 : std_logic := '0';
  signal q9 : std_logic := '0';
  signal qdrive : std_logic := '0';
  signal qs0 : std_logic := '0';
  signal qs1 : std_logic := '0';
  signal r0 : std_logic := '0';
  signal r1 : std_logic := '0';
  signal r10 : std_logic := '0';
  signal r11 : std_logic := '0';
  signal r12 : std_logic := '0';
  signal r13 : std_logic := '0';
  signal r14 : std_logic := '0';
  signal r15 : std_logic := '0';
  signal r16 : std_logic := '0';
  signal r17 : std_logic := '0';
  signal r18 : std_logic := '0';
  signal r19 : std_logic := '0';
  signal r2 : std_logic := '0';
  signal r20 : std_logic := '0';
  signal r21 : std_logic := '0';
  signal r22 : std_logic := '0';
  signal r23 : std_logic := '0';
  signal r24 : std_logic := '0';
  signal r25 : std_logic := '0';
  signal r26 : std_logic := '0';
  signal r27 : std_logic := '0';
  signal r28 : std_logic := '0';
  signal r29 : std_logic := '0';
  signal r3 : std_logic := '0';
  signal r30 : std_logic := '0';
  signal r31 : std_logic := '0';
  signal r4 : std_logic := '0';
  signal r5 : std_logic := '0';
  signal r6 : std_logic := '0';
  signal r7 : std_logic := '0';
  signal r8 : std_logic := '0';
  signal r9 : std_logic := '0';
  signal ramdisable : std_logic := '0';
  signal rdcyc : std_logic := '0';
  signal reset : std_logic := '0';
  signal reta0 : std_logic := '0';
  signal reta1 : std_logic := '0';
  signal reta10 : std_logic := '0';
  signal reta11 : std_logic := '0';
  signal reta12 : std_logic := '0';
  signal reta13 : std_logic := '0';
  signal reta2 : std_logic := '0';
  signal reta3 : std_logic := '0';
  signal reta4 : std_logic := '0';
  signal reta5 : std_logic := '0';
  signal reta6 : std_logic := '0';
  signal reta7 : std_logic := '0';
  signal reta8 : std_logic := '0';
  signal reta9 : std_logic := '0';
  signal run : std_logic := '0';
  signal s0 : std_logic := '0';
  signal s1 : std_logic := '0';
  signal s2a : std_logic := '0';
  signal s2b : std_logic := '0';
  signal s3a : std_logic := '0';
  signal s3b : std_logic := '0';
  signal s4 : std_logic := '0';
  signal sa0 : std_logic := '0';
  signal sa1 : std_logic := '0';
  signal sa10 : std_logic := '0';
  signal sa11 : std_logic := '0';
  signal sa12 : std_logic := '0';
  signal sa13 : std_logic := '0';
  signal sa14 : std_logic := '0';
  signal sa15 : std_logic := '0';
  signal sa16 : std_logic := '0';
  signal sa17 : std_logic := '0';
  signal sa18 : std_logic := '0';
  signal sa19 : std_logic := '0';
  signal sa2 : std_logic := '0';
  signal sa20 : std_logic := '0';
  signal sa21 : std_logic := '0';
  signal sa22 : std_logic := '0';
  signal sa23 : std_logic := '0';
  signal sa24 : std_logic := '0';
  signal sa25 : std_logic := '0';
  signal sa26 : std_logic := '0';
  signal sa27 : std_logic := '0';
  signal sa28 : std_logic := '0';
  signal sa29 : std_logic := '0';
  signal sa3 : std_logic := '0';
  signal sa30 : std_logic := '0';
  signal sa31 : std_logic := '0';
  signal sa4 : std_logic := '0';
  signal sa5 : std_logic := '0';
  signal sa6 : std_logic := '0';
  signal sa7 : std_logic := '0';
  signal sa8 : std_logic := '0';
  signal sa9 : std_logic := '0';
  signal sint : std_logic := '0';
  signal sintr : std_logic := '0';
  signal spc0 : std_logic := '0';
  signal spc1 : std_logic := '0';
  signal spc10 : std_logic := '0';
  signal spc11 : std_logic := '0';
  signal spc12 : std_logic := '0';
  signal spc13 : std_logic := '0';
  signal spc14 : std_logic := '0';
  signal spc15 : std_logic := '0';
  signal spc16 : std_logic := '0';
  signal spc17 : std_logic := '0';
  signal spc18 : std_logic := '0';
  signal spc1a : std_logic := '0';
  signal spc2 : std_logic := '0';
  signal spc3 : std_logic := '0';
  signal spc4 : std_logic := '0';
  signal spc5 : std_logic := '0';
  signal spc6 : std_logic := '0';
  signal spc7 : std_logic := '0';
  signal spc8 : std_logic := '0';
  signal spc9 : std_logic := '0';
  signal spcdrive : std_logic := '0';
  signal spcenb : std_logic := '0';
  signal spcmung : std_logic := '0';
  signal spco0 : std_logic := '0';
  signal spco1 : std_logic := '0';
  signal spco10 : std_logic := '0';
  signal spco11 : std_logic := '0';
  signal spco12 : std_logic := '0';
  signal spco13 : std_logic := '0';
  signal spco14 : std_logic := '0';
  signal spco15 : std_logic := '0';
  signal spco16 : std_logic := '0';
  signal spco17 : std_logic := '0';
  signal spco18 : std_logic := '0';
  signal spco2 : std_logic := '0';
  signal spco3 : std_logic := '0';
  signal spco4 : std_logic := '0';
  signal spco5 : std_logic := '0';
  signal spco6 : std_logic := '0';
  signal spco7 : std_logic := '0';
  signal spco8 : std_logic := '0';
  signal spco9 : std_logic := '0';
  signal spcopar : std_logic := '0';
  signal spcpar : std_logic := '0';
  signal spcparh : std_logic := '0';
  signal spcparok : std_logic := '0';
  signal spcptr0 : std_logic := '0';
  signal spcptr1 : std_logic := '0';
  signal spcptr2 : std_logic := '0';
  signal spcptr3 : std_logic := '0';
  signal spcptr4 : std_logic := '0';
  signal spcw0 : std_logic := '0';
  signal spcw1 : std_logic := '0';
  signal spcw10 : std_logic := '0';
  signal spcw11 : std_logic := '0';
  signal spcw12 : std_logic := '0';
  signal spcw13 : std_logic := '0';
  signal spcw14 : std_logic := '0';
  signal spcw15 : std_logic := '0';
  signal spcw16 : std_logic := '0';
  signal spcw17 : std_logic := '0';
  signal spcw18 : std_logic := '0';
  signal spcw2 : std_logic := '0';
  signal spcw3 : std_logic := '0';
  signal spcw4 : std_logic := '0';
  signal spcw5 : std_logic := '0';
  signal spcw6 : std_logic := '0';
  signal spcw7 : std_logic := '0';
  signal spcw8 : std_logic := '0';
  signal spcw9 : std_logic := '0';
  signal spcwpar : std_logic := '0';
  signal spcwparh : std_logic := '0';
  signal spcwpass : std_logic := '0';
  signal speed0 : std_logic := '0';
  signal speed0a : std_logic := '0';
  signal speed1 : std_logic := '0';
  signal speed1a : std_logic := '0';
  signal speedclk : std_logic := '0';
  signal spush : std_logic := '0';
  signal spushd : std_logic := '0';
  signal spy0 : std_logic := '0';
  signal spy1 : std_logic := '0';
  signal spy10 : std_logic := '0';
  signal spy11 : std_logic := '0';
  signal spy12 : std_logic := '0';
  signal spy13 : std_logic := '0';
  signal spy14 : std_logic := '0';
  signal spy15 : std_logic := '0';
  signal spy2 : std_logic := '0';
  signal spy3 : std_logic := '0';
  signal spy4 : std_logic := '0';
  signal spy5 : std_logic := '0';
  signal spy6 : std_logic := '0';
  signal spy7 : std_logic := '0';
  signal spy8 : std_logic := '0';
  signal spy9 : std_logic := '0';
  signal srclc : std_logic := '0';
  signal srcm : std_logic := '0';
  signal srcmap : std_logic := '0';
  signal srcmd : std_logic := '0';
  signal srcpdlidx : std_logic := '0';
  signal srcpdlptr : std_logic := '0';
  signal srcq : std_logic := '0';
  signal srcvma : std_logic := '0';
  signal srun : std_logic := '0';
  signal ssdone : std_logic := '0';
  signal sspeed0 : std_logic := '0';
  signal sspeed1 : std_logic := '0';
  signal sstep : std_logic := '0';
  signal st0 : std_logic := '0';
  signal st1 : std_logic := '0';
  signal st10 : std_logic := '0';
  signal st11 : std_logic := '0';
  signal st12 : std_logic := '0';
  signal st13 : std_logic := '0';
  signal st14 : std_logic := '0';
  signal st15 : std_logic := '0';
  signal st16 : std_logic := '0';
  signal st17 : std_logic := '0';
  signal st18 : std_logic := '0';
  signal st19 : std_logic := '0';
  signal st2 : std_logic := '0';
  signal st20 : std_logic := '0';
  signal st21 : std_logic := '0';
  signal st22 : std_logic := '0';
  signal st23 : std_logic := '0';
  signal st24 : std_logic := '0';
  signal st25 : std_logic := '0';
  signal st26 : std_logic := '0';
  signal st27 : std_logic := '0';
  signal st28 : std_logic := '0';
  signal st29 : std_logic := '0';
  signal st3 : std_logic := '0';
  signal st30 : std_logic := '0';
  signal st31 : std_logic := '0';
  signal st4 : std_logic := '0';
  signal st5 : std_logic := '0';
  signal st6 : std_logic := '0';
  signal st7 : std_logic := '0';
  signal st8 : std_logic := '0';
  signal st9 : std_logic := '0';
  signal stathenb : std_logic := '0';
  signal statstop : std_logic := '0';
  signal step : std_logic := '0';
  signal tilt0 : std_logic := '0';
  signal tilt1 : std_logic := '0';
  signal tpclk : std_logic := '0';
  signal tprend : std_logic := '0';
  signal tptse : std_logic := '0';
  signal tpwp : std_logic := '0';
  signal tpwpiram : std_logic := '0';
  signal trapa : std_logic := '0';
  signal trapb : std_logic := '0';
  signal trapenb : std_logic := '0';
  signal tse1a : std_logic := '0';
  signal tse1b : std_logic := '0';
  signal tse2 : std_logic := '0';
  signal tse3a : std_logic := '0';
  signal tse4a : std_logic := '0';
  signal tse4b : std_logic := '0';
  signal v0parok : std_logic := '0';
  signal vm0pari : std_logic := '0';
  signal vm1mpar : std_logic := '0';
  signal vm1pari : std_logic := '0';
  signal vmap0a : std_logic := '0';
  signal vmap0b : std_logic := '0';
  signal vmap1a : std_logic := '0';
  signal vmap1b : std_logic := '0';
  signal vmap2a : std_logic := '0';
  signal vmap2b : std_logic := '0';
  signal vmap3a : std_logic := '0';
  signal vmap3b : std_logic := '0';
  signal vmap4a : std_logic := '0';
  signal vmap4b : std_logic := '0';
  signal vmasela : std_logic := '0';
  signal vmaselb : std_logic := '0';
  signal vmo18 : std_logic := '0';
  signal vmo19 : std_logic := '0';
  signal vmopar : std_logic := '0';
  signal vmoparck : std_logic := '0';
  signal vmoparl : std_logic := '0';
  signal vmoparm : std_logic := '0';
  signal vmoparodd : std_logic := '0';
  signal vmoparok : std_logic := '0';
  signal vpari : std_logic := '0';
  signal wadr0 : std_logic := '0';
  signal wadr1 : std_logic := '0';
  signal wadr2 : std_logic := '0';
  signal wadr3 : std_logic := '0';
  signal wadr4 : std_logic := '0';
  signal wadr5 : std_logic := '0';
  signal wadr6 : std_logic := '0';
  signal wadr7 : std_logic := '0';
  signal wadr8 : std_logic := '0';
  signal wadr9 : std_logic := '0';
  signal wmap : std_logic := '0';
  signal wmapd : std_logic := '0';
  signal wp1a : std_logic := '0';
  signal wp1b : std_logic := '0';
  signal wp2 : std_logic := '0';
  signal wp3a : std_logic := '0';
  signal wp4a : std_logic := '0';
  signal wp4b : std_logic := '0';
  signal wp4c : std_logic := '0';
  signal wp5a : std_logic := '0';
  signal wp5b : std_logic := '0';
  signal wp5c : std_logic := '0';
  signal wp5d : std_logic := '0';
  signal wpc0 : std_logic := '0';
  signal wpc1 : std_logic := '0';
  signal wpc10 : std_logic := '0';
  signal wpc11 : std_logic := '0';
  signal wpc12 : std_logic := '0';
  signal wpc13 : std_logic := '0';
  signal wpc2 : std_logic := '0';
  signal wpc3 : std_logic := '0';
  signal wpc4 : std_logic := '0';
  signal wpc5 : std_logic := '0';
  signal wpc6 : std_logic := '0';
  signal wpc7 : std_logic := '0';
  signal wpc8 : std_logic := '0';
  signal wpc9 : std_logic := '0';
  signal wrcyc : std_logic := '0';
  signal xout11 : std_logic := '0';
  signal xout15 : std_logic := '0';
  signal xout19 : std_logic := '0';
  signal xout23 : std_logic := '0';
  signal xout27 : std_logic := '0';
  signal xout3 : std_logic := '0';
  signal xout31 : std_logic := '0';
  signal xout7 : std_logic := '0';
  signal xx0 : std_logic := '0';
  signal xx1 : std_logic := '0';
  signal yout11 : std_logic := '0';
  signal yout15 : std_logic := '0';
  signal yout19 : std_logic := '0';
  signal yout23 : std_logic := '0';
  signal yout27 : std_logic := '0';
  signal yout3 : std_logic := '0';
  signal yout31 : std_logic := '0';
  signal yout7 : std_logic := '0';
  signal yy0 : std_logic := '0';
  signal yy1 : std_logic := '0';
  signal zero16 : std_logic := '0';
begin

--- Clock Generation (clkgen)
  i_clock1 : entity icmem_book.clock1(ttl) port map(\-clock_reset_b\ => \-clock_reset_b\, \-tpdone\ => \-tpdone\, \-hang\ => \-hang\, cyclecompleted => cyclecompleted, \-tpr0\ => \-tpr0\, \-tpr40\ => \-tpr40\, gnd => gnd, \-tprend\ => \-tprend\, \-tpw20\ => \-tpw20\, \-tpw40\ => \-tpw40\, \-tpw50\ => \-tpw50\, \-tpw30\ => \-tpw30\, \-tpw10\ => \-tpw10\, \-tpw60\ => \-tpw60\, \-tpw70\ => \-tpw70\, \-tpw75\ => \-tpw75\, \-tpw65\ => \-tpw65\, \-tpw55\ => \-tpw55\, \-tpw30a\ => \-tpw30a\, \-tpw40a\ => \-tpw40a\, \-tpw45\ => \-tpw45\, \-tpw35\ => \-tpw35\, \-tpw25\ => \-tpw25\, \-tpr100\ => \-tpr100\, \-tpr140\ => \-tpr140\, \-tpr160\ => \-tpr160\, tprend => tprend, sspeed1 => sspeed1, sspeed0 => sspeed0, \-ilong\ => \-ilong\, \-tpr75\ => \-tpr75\, \-tpr115\ => \-tpr115\, \-tpr85\ => \-tpr85\, \-tpr125\ => \-tpr125\, \-tpr10\ => \-tpr10\, \-tpr20a\ => \-tpr20a\, \-tpr25\ => \-tpr25\, \-tpr15\ => \-tpr15\, \-tpr5\ => \-tpr5\, \-tpr80\ => \-tpr80\, \-tpr60\ => \-tpr60\, \-tpr20\ => \-tpr20\, \-tpr180\ => \-tpr180\, \-tpr200\ => \-tpr200\, \-tpr120\ => \-tpr120\, \-tpr110\ => \-tpr110\, \-tpr120a\ => \-tpr120a\, \-tpr105\ => \-tpr105\, \-tpr70\ => \-tpr70\, \-tpr80a\ => \-tpr80a\, \-tpr65\ => \-tpr65\);
  i_clock2 : entity icmem_book.clock2(ttl) port map(clk4 => clk4, \-clk0\ => \-clk0\, gnd => gnd, mclk7 => mclk7, \-mclk0\ => \-mclk0\, \-wp1\ => \-wp1\, tpwp => tpwp, \-wp2\ => \-wp2\, \-wp3\ => \-wp3\, \-wp4\ => \-wp4\, \-tprend\ => \-tprend\, tpclk => tpclk, \-tptse\ => \-tptse\, \-tpr25\ => \-tpr25\, \-clock_reset_b\ => \-clock_reset_b\, tptse => tptse, \-tpw70\ => \-tpw70\, \-tpclk\ => \-tpclk\, \-tpr0\ => \-tpr0\, \-tpr5\ => \-tpr5\, \-tpw30\ => \-tpw30\, \machruna_l\ => \machruna_l\, tpwpiram => tpwpiram, \-wp5\ => \-wp5\, clk5 => clk5, mclk5 => mclk5, \-tpw45\ => \-tpw45\, \-tse1\ => \-tse1\, \-tse2\ => \-tse2\, \-tse3\ => \-tse3\, \-tse4\ => \-tse4\, clk1 => clk1, clk2 => clk2, clk3 => clk3, mclk1 => mclk1, machrun => machrun, hi1 => hi1);
  i_clockd : entity cadr_book.clockd(ttl) port map(\-clk1\ => \-clk1\, hi12 => hi12, clk1a => clk1a, reset => reset, \-reset\ => \-reset\, mclk1a => mclk1a, \-mclk1\ => \-mclk1\, mclk1 => mclk1, clk1 => clk1, \-wp1\ => \-wp1\, wp1b => wp1b, wp1a => wp1a, tse1b => tse1b, \-tse1\ => \-tse1\, tse1a => tse1a, hi1 => hi1, hi2 => hi2, hi3 => hi3, hi4 => hi4, hi5 => hi5, hi6 => hi6, hi7 => hi7, \-upperhighok\ => \-upperhighok\, hi8 => hi8, hi9 => hi9, hi10 => hi10, hi11 => hi11, lcry3 => lcry3, \-lcry3\ => \-lcry3\, clk2 => clk2, \-clk2c\ => \-clk2c\, \-clk2a\ => \-clk2a\, wp2 => wp2, \-wp2\ => \-wp2\, tse2 => tse2, \-tse2\ => \-tse2\, clk2a => clk2a, clk2b => clk2b, clk2c => clk2c, \-clk3a\ => \-clk3a\, clk3a => clk3a, clk3b => clk3b, clk3c => clk3c, clk3 => clk3, \-clk3g\ => \-clk3g\, \-clk3d\ => \-clk3d\, wp3a => wp3a, \-wp3\ => \-wp3\, tse3a => tse3a, \-tse3\ => \-tse3\, clk3d => clk3d, clk3e => clk3e, clk3f => clk3f, \-clk4a\ => \-clk4a\, clk4a => clk4a, clk4b => clk4b, clk4c => clk4c, clk4 => clk4, \-clk4e\ => \-clk4e\, \-clk4d\ => \-clk4d\, wp4c => wp4c, \-wp4\ => \-wp4\, wp4b => wp4b, wp4a => wp4a, clk4d => clk4d, clk4e => clk4e, clk4f => clk4f, \-tse4\ => \-tse4\, tse4b => tse4b, tse4a => tse4a, srcpdlptr => srcpdlptr, \-srcpdlptr\ => \-srcpdlptr\, srcpdlidx => srcpdlidx, \-srcpdlidx\ => \-srcpdlidx\);


--- Microinstruction Fetch (imem?)
  i_ictl : entity icmem_book.ictl(ttl) port map(ramdisable => ramdisable, hi1 => hi1, \-iwriteda\ => \-iwriteda\, \-promdisabled\ => \-promdisabled\, idebug => idebug, iwriteda => iwriteda, promdisabled => promdisabled, \-wp5\ => \-wp5\, wp5d => wp5d, wp5c => wp5c, wp5b => wp5b, wp5a => wp5a, pc0 => pc0, \-pcb0\ => \-pcb0\, pc1 => pc1, \-pcb1\ => \-pcb1\, pc2 => pc2, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, pc3 => pc3, \-pcb4\ => \-pcb4\, pc4 => pc4, \-pcb5\ => \-pcb5\, pc5 => pc5, \-iwea\ => \-iwea\, \-iweb\ => \-iweb\, \-iwei\ => \-iwei\, \-iwej\ => \-iwej\, pc13 => pc13, \-pc13b\ => \-pc13b\, pc12 => pc12, \-pc12b\ => \-pc12b\, \-iwrited\ => \-iwrited\, iwritedd => iwritedd, iwritedc => iwritedc, iwritedb => iwritedb, pc6 => pc6, \-pcb6\ => \-pcb6\, pc7 => pc7, \-pcb7\ => \-pcb7\, pc8 => pc8, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, pc9 => pc9, \-pcb10\ => \-pcb10\, pc10 => pc10, \-pcb11\ => \-pcb11\, pc11 => pc11, \-ice3a\ => \-ice3a\, \-ice2a\ => \-ice2a\, \-ice1a\ => \-ice1a\, \-ice0a\ => \-ice0a\, \-ice0b\ => \-ice0b\, \-ice1b\ => \-ice1b\, \-ice2b\ => \-ice2b\, \-ice3b\ => \-ice3b\, \-iwec\ => \-iwec\, \-iwed\ => \-iwed\, \-iwek\ => \-iwek\, \-iwel\ => \-iwel\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-iwee\ => \-iwee\, \-iwef\ => \-iwef\, \-iwem\ => \-iwem\, \-iwen\ => \-iwen\, \-ice3c\ => \-ice3c\, \-ice2c\ => \-ice2c\, \-ice1c\ => \-ice1c\, \-ice0c\ => \-ice0c\, \-ice0d\ => \-ice0d\, \-ice1d\ => \-ice1d\, \-ice2d\ => \-ice2d\, \-ice3d\ => \-ice3d\, \-iweg\ => \-iweg\, \-iweh\ => \-iweh\, \-iweo\ => \-iweo\, \-iwep\ => \-iwep\);
  i_iram00 : entity icmem_book.iram00(ttl) port map(pc0a => pc0a, pc1a => pc1a, pc2a => pc2a, pc3a => pc3a, pc4a => pc4a, pc5a => pc5a, i10 => i10, \-iwea\ => \-iwea\, \-ice0a\ => \-ice0a\, iwr10 => iwr10, pc11a => pc11a, pc10a => pc10a, pc9a => pc9a, pc8a => pc8a, pc7a => pc7a, pc6a => pc6a, i11 => i11, iwr11 => iwr11, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i5 => i5, iwr5 => iwr5, i6 => i6, iwr6 => iwr6, i7 => i7, iwr7 => iwr7, i8 => i8, iwr8 => iwr8, i9 => i9, iwr9 => iwr9, i0 => i0, iwr0 => iwr0, i1 => i1, iwr1 => iwr1, i2 => i2, iwr2 => iwr2, i3 => i3, iwr3 => iwr3, i4 => i4, iwr4 => iwr4);
  i_iram01 : entity icmem_book.iram01(ttl) port map(pc0b => pc0b, pc1b => pc1b, pc2b => pc2b, pc3b => pc3b, pc4b => pc4b, pc5b => pc5b, i10 => i10, \-iweb\ => \-iweb\, \-ice1a\ => \-ice1a\, iwr10 => iwr10, pc11b => pc11b, pc10b => pc10b, pc9b => pc9b, pc8b => pc8b, pc7b => pc7b, pc6b => pc6b, i11 => i11, iwr11 => iwr11, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i5 => i5, iwr5 => iwr5, i6 => i6, iwr6 => iwr6, i7 => i7, iwr7 => iwr7, i8 => i8, iwr8 => iwr8, i9 => i9, iwr9 => iwr9, i0 => i0, iwr0 => iwr0, i1 => i1, iwr1 => iwr1, i2 => i2, iwr2 => iwr2, i3 => i3, iwr3 => iwr3, i4 => i4, iwr4 => iwr4);
  i_iram02 : entity icmem_book.iram02(ttl) port map(pc0c => pc0c, pc1c => pc1c, pc2c => pc2c, pc3c => pc3c, pc4c => pc4c, pc5c => pc5c, i10 => i10, \-iwec\ => \-iwec\, \-ice2a\ => \-ice2a\, iwr10 => iwr10, pc11c => pc11c, pc10c => pc10c, pc9c => pc9c, pc8c => pc8c, pc7c => pc7c, pc6c => pc6c, i11 => i11, iwr11 => iwr11, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i5 => i5, iwr5 => iwr5, i6 => i6, iwr6 => iwr6, i7 => i7, iwr7 => iwr7, i8 => i8, iwr8 => iwr8, i9 => i9, iwr9 => iwr9, i0 => i0, iwr0 => iwr0, i1 => i1, iwr1 => iwr1, i2 => i2, iwr2 => iwr2, i3 => i3, iwr3 => iwr3, i4 => i4, iwr4 => iwr4);
  i_iram03 : entity icmem_book.iram03(ttl) port map(pc0d => pc0d, pc1d => pc1d, pc2d => pc2d, pc3d => pc3d, pc4d => pc4d, pc5d => pc5d, i10 => i10, \-iwed\ => \-iwed\, \-ice3a\ => \-ice3a\, iwr10 => iwr10, pc11d => pc11d, pc10d => pc10d, pc9d => pc9d, pc8d => pc8d, pc7d => pc7d, pc6d => pc6d, i11 => i11, iwr11 => iwr11, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i5 => i5, iwr5 => iwr5, i6 => i6, iwr6 => iwr6, i7 => i7, iwr7 => iwr7, i8 => i8, iwr8 => iwr8, i9 => i9, iwr9 => iwr9, i0 => i0, iwr0 => iwr0, i1 => i1, iwr1 => iwr1, i2 => i2, iwr2 => iwr2, i3 => i3, iwr3 => iwr3, i4 => i4, iwr4 => iwr4);
  i_iram10 : entity icmem_book.iram10(ttl) port map(pc0e => pc0e, pc1e => pc1e, pc2e => pc2e, pc3e => pc3e, pc4e => pc4e, pc5e => pc5e, i22 => i22, \-iwee\ => \-iwee\, \-ice0b\ => \-ice0b\, iwr22 => iwr22, pc11e => pc11e, pc10e => pc10e, pc9e => pc9e, pc8e => pc8e, pc7e => pc7e, pc6e => pc6e, i23 => i23, iwr23 => iwr23, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i17 => i17, iwr17 => iwr17, i18 => i18, iwr18 => iwr18, i19 => i19, iwr19 => iwr19, i20 => i20, iwr20 => iwr20, i21 => i21, iwr21 => iwr21, i12 => i12, iwr12 => iwr12, i13 => i13, iwr13 => iwr13, i14 => i14, iwr14 => iwr14, i15 => i15, iwr15 => iwr15, i16 => i16, iwr16 => iwr16);
  i_iram11 : entity icmem_book.iram11(ttl) port map(pc0f => pc0f, pc1f => pc1f, pc2f => pc2f, pc3f => pc3f, pc4f => pc4f, pc5f => pc5f, i22 => i22, \-iwef\ => \-iwef\, \-ice1b\ => \-ice1b\, iwr22 => iwr22, pc11f => pc11f, pc10f => pc10f, pc9f => pc9f, pc8f => pc8f, pc7f => pc7f, pc6f => pc6f, i23 => i23, iwr23 => iwr23, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i17 => i17, iwr17 => iwr17, i18 => i18, iwr18 => iwr18, i19 => i19, iwr19 => iwr19, i20 => i20, iwr20 => iwr20, i21 => i21, iwr21 => iwr21, i12 => i12, iwr12 => iwr12, i13 => i13, iwr13 => iwr13, i14 => i14, iwr14 => iwr14, i15 => i15, iwr15 => iwr15, i16 => i16, iwr16 => iwr16);
  i_iram12 : entity icmem_book.iram12(ttl) port map(pc0g => pc0g, pc1g => pc1g, pc2g => pc2g, pc3g => pc3g, pc4g => pc4g, pc5g => pc5g, i22 => i22, \-iweg\ => \-iweg\, \-ice2b\ => \-ice2b\, iwr22 => iwr22, pc11g => pc11g, pc10g => pc10g, pc9g => pc9g, pc8g => pc8g, pc7g => pc7g, pc6g => pc6g, i23 => i23, iwr23 => iwr23, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i17 => i17, iwr17 => iwr17, i18 => i18, iwr18 => iwr18, i19 => i19, iwr19 => iwr19, i20 => i20, iwr20 => iwr20, i21 => i21, iwr21 => iwr21, i12 => i12, iwr12 => iwr12, i13 => i13, iwr13 => iwr13, i14 => i14, iwr14 => iwr14, i15 => i15, iwr15 => iwr15, i16 => i16, iwr16 => iwr16);
  i_iram13 : entity icmem_book.iram13(ttl) port map(pc0h => pc0h, pc1h => pc1h, pc2h => pc2h, pc3h => pc3h, pc4h => pc4h, pc5h => pc5h, i22 => i22, \-iweh\ => \-iweh\, \-ice3b\ => \-ice3b\, iwr22 => iwr22, pc11h => pc11h, pc10h => pc10h, pc9h => pc9h, pc8h => pc8h, pc7h => pc7h, pc6h => pc6h, i23 => i23, iwr23 => iwr23, \-pcb6\ => \-pcb6\, \-pcb7\ => \-pcb7\, \-pcb8\ => \-pcb8\, \-pcb9\ => \-pcb9\, \-pcb10\ => \-pcb10\, \-pcb11\ => \-pcb11\, \-pcb0\ => \-pcb0\, \-pcb1\ => \-pcb1\, \-pcb2\ => \-pcb2\, \-pcb3\ => \-pcb3\, \-pcb4\ => \-pcb4\, \-pcb5\ => \-pcb5\, i17 => i17, iwr17 => iwr17, i18 => i18, iwr18 => iwr18, i19 => i19, iwr19 => iwr19, i20 => i20, iwr20 => iwr20, i21 => i21, iwr21 => iwr21, i12 => i12, iwr12 => iwr12, i13 => i13, iwr13 => iwr13, i14 => i14, iwr14 => iwr14, i15 => i15, iwr15 => iwr15, i16 => i16, iwr16 => iwr16);
  i_iram20 : entity icmem_book.iram20(ttl) port map(pc0i => pc0i, pc1i => pc1i, pc2i => pc2i, pc3i => pc3i, pc4i => pc4i, pc5i => pc5i, i31 => i31, \-iwei\ => \-iwei\, \-ice0c\ => \-ice0c\, iwr31 => iwr31, pc11i => pc11i, pc10i => pc10i, pc9i => pc9i, pc8i => pc8i, pc7i => pc7i, pc6i => pc6i, i32 => i32, iwr32 => iwr32, i33 => i33, iwr33 => iwr33, i34 => i34, iwr34 => iwr34, i35 => i35, iwr35 => iwr35, i26 => i26, iwr26 => iwr26, i27 => i27, iwr27 => iwr27, i28 => i28, iwr28 => iwr28, i29 => i29, iwr29 => iwr29, i30 => i30, iwr30 => iwr30, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i24 => i24, iwr24 => iwr24, i25 => i25, iwr25 => iwr25);
  i_iram21 : entity icmem_book.iram21(ttl) port map(pc0j => pc0j, pc1j => pc1j, pc2j => pc2j, pc3j => pc3j, pc4j => pc4j, pc5j => pc5j, i31 => i31, \-iwej\ => \-iwej\, \-ice1c\ => \-ice1c\, iwr31 => iwr31, pc11j => pc11j, pc10j => pc10j, pc9j => pc9j, pc8j => pc8j, pc7j => pc7j, pc6j => pc6j, i32 => i32, iwr32 => iwr32, i33 => i33, iwr33 => iwr33, i34 => i34, iwr34 => iwr34, i35 => i35, iwr35 => iwr35, i26 => i26, iwr26 => iwr26, i27 => i27, iwr27 => iwr27, i28 => i28, iwr28 => iwr28, i29 => i29, iwr29 => iwr29, i30 => i30, iwr30 => iwr30, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i24 => i24, iwr24 => iwr24, i25 => i25, iwr25 => iwr25);
  i_iram22 : entity icmem_book.iram22(ttl) port map(pc0k => pc0k, pc1k => pc1k, pc2k => pc2k, pc3k => pc3k, pc4k => pc4k, pc5k => pc5k, i31 => i31, \-iwek\ => \-iwek\, \-ice2c\ => \-ice2c\, iwr31 => iwr31, pc11k => pc11k, pc10k => pc10k, pc9k => pc9k, pc8k => pc8k, pc7k => pc7k, pc6k => pc6k, i32 => i32, iwr32 => iwr32, i33 => i33, iwr33 => iwr33, i34 => i34, iwr34 => iwr34, i35 => i35, iwr35 => iwr35, i26 => i26, iwr26 => iwr26, i27 => i27, iwr27 => iwr27, i28 => i28, iwr28 => iwr28, i29 => i29, iwr29 => iwr29, i30 => i30, iwr30 => iwr30, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i24 => i24, iwr24 => iwr24, i25 => i25, iwr25 => iwr25);
  i_iram23 : entity icmem_book.iram23(ttl) port map(pc0l => pc0l, pc1l => pc1l, pc2l => pc2l, pc3l => pc3l, pc4l => pc4l, pc5l => pc5l, i31 => i31, \-iwel\ => \-iwel\, \-ice3c\ => \-ice3c\, iwr31 => iwr31, pc11l => pc11l, pc10l => pc10l, pc9l => pc9l, pc8l => pc8l, pc7l => pc7l, pc6l => pc6l, i32 => i32, iwr32 => iwr32, i33 => i33, iwr33 => iwr33, i34 => i34, iwr34 => iwr34, i35 => i35, iwr35 => iwr35, i26 => i26, iwr26 => iwr26, i27 => i27, iwr27 => iwr27, i28 => i28, iwr28 => iwr28, i29 => i29, iwr29 => iwr29, i30 => i30, iwr30 => iwr30, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i24 => i24, iwr24 => iwr24, i25 => i25, iwr25 => iwr25);
  i_iram30 : entity icmem_book.iram30(ttl) port map(pc0m => pc0m, pc1m => pc1m, pc2m => pc2m, pc3m => pc3m, pc4m => pc4m, pc5m => pc5m, i44 => i44, \-iwem\ => \-iwem\, \-ice0d\ => \-ice0d\, iwr44 => iwr44, pc11m => pc11m, pc10m => pc10m, pc9m => pc9m, pc8m => pc8m, pc7m => pc7m, pc6m => pc6m, i45 => i45, iwr45 => iwr45, i46 => i46, iwr46 => iwr46, i47 => i47, iwr47 => iwr47, i48 => i48, iwr48 => iwr48, i39 => i39, iwr39 => iwr39, i40 => i40, iwr40 => iwr40, i41 => i41, iwr41 => iwr41, i42 => i42, iwr42 => iwr42, i43 => i43, iwr43 => iwr43, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i36 => i36, iwr36 => iwr36, i37 => i37, iwr37 => iwr37, i38 => i38, iwr38 => iwr38);
  i_iram31 : entity icmem_book.iram31(ttl) port map(pc0n => pc0n, pc1n => pc1n, pc2n => pc2n, pc3n => pc3n, pc4n => pc4n, pc5n => pc5n, i44 => i44, \-iwen\ => \-iwen\, \-ice1d\ => \-ice1d\, iwr44 => iwr44, pc11n => pc11n, pc10n => pc10n, pc9n => pc9n, pc8n => pc8n, pc7n => pc7n, pc6n => pc6n, i45 => i45, iwr45 => iwr45, i46 => i46, iwr46 => iwr46, i47 => i47, iwr47 => iwr47, i48 => i48, iwr48 => iwr48, i39 => i39, iwr39 => iwr39, i40 => i40, iwr40 => iwr40, i41 => i41, iwr41 => iwr41, i42 => i42, iwr42 => iwr42, i43 => i43, iwr43 => iwr43, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i36 => i36, iwr36 => iwr36, i37 => i37, iwr37 => iwr37, i38 => i38, iwr38 => iwr38);
  i_iram32 : entity icmem_book.iram32(ttl) port map(pc0o => pc0o, pc1o => pc1o, pc2o => pc2o, pc3o => pc3o, pc4o => pc4o, pc5o => pc5o, i44 => i44, \-iweo\ => \-iweo\, \-ice2d\ => \-ice2d\, iwr44 => iwr44, pc11o => pc11o, pc10o => pc10o, pc9o => pc9o, pc8o => pc8o, pc7o => pc7o, pc6o => pc6o, i45 => i45, iwr45 => iwr45, i46 => i46, iwr46 => iwr46, i47 => i47, iwr47 => iwr47, i48 => i48, iwr48 => iwr48, i39 => i39, iwr39 => iwr39, i40 => i40, iwr40 => iwr40, i41 => i41, iwr41 => iwr41, i42 => i42, iwr42 => iwr42, i43 => i43, iwr43 => iwr43, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i36 => i36, iwr36 => iwr36, i37 => i37, iwr37 => iwr37, i38 => i38, iwr38 => iwr38);
  i_iram33 : entity icmem_book.iram33(ttl) port map(pc0p => pc0p, pc1p => pc1p, pc2p => pc2p, pc3p => pc3p, pc4p => pc4p, pc5p => pc5p, i44 => i44, \-iwep\ => \-iwep\, \-ice3d\ => \-ice3d\, iwr44 => iwr44, pc11p => pc11p, pc10p => pc10p, pc9p => pc9p, pc8p => pc8p, pc7p => pc7p, pc6p => pc6p, i45 => i45, iwr45 => iwr45, i46 => i46, iwr46 => iwr46, i47 => i47, iwr47 => iwr47, i48 => i48, iwr48 => iwr48, i39 => i39, iwr39 => iwr39, i40 => i40, iwr40 => iwr40, i41 => i41, iwr41 => iwr41, i42 => i42, iwr42 => iwr42, i43 => i43, iwr43 => iwr43, \-pcc6\ => \-pcc6\, \-pcc7\ => \-pcc7\, \-pcc8\ => \-pcc8\, \-pcc9\ => \-pcc9\, \-pcc10\ => \-pcc10\, \-pcc11\ => \-pcc11\, \-pcc0\ => \-pcc0\, \-pcc1\ => \-pcc1\, \-pcc2\ => \-pcc2\, \-pcc3\ => \-pcc3\, \-pcc4\ => \-pcc4\, \-pcc5\ => \-pcc5\, i36 => i36, iwr36 => iwr36, i37 => i37, iwr37 => iwr37, i38 => i38, iwr38 => iwr38);
  i_iwr : entity cadr_book.iwr(ttl) port map(gnd => gnd, iwr47 => iwr47, aa15 => aa15, aa14 => aa14, iwr46 => iwr46, iwr45 => iwr45, aa13 => aa13, aa12 => aa12, iwr44 => iwr44, clk2c => clk2c, iwr43 => iwr43, aa11 => aa11, aa10 => aa10, iwr42 => iwr42, iwr41 => iwr41, aa9 => aa9, aa8 => aa8, iwr40 => iwr40, iwr39 => iwr39, aa7 => aa7, aa6 => aa6, iwr38 => iwr38, iwr37 => iwr37, aa5 => aa5, aa4 => aa4, iwr36 => iwr36, iwr35 => iwr35, aa3 => aa3, aa2 => aa2, iwr34 => iwr34, iwr33 => iwr33, aa1 => aa1, aa0 => aa0, iwr32 => iwr32, iwr15 => iwr15, m15 => m15, m14 => m14, iwr14 => iwr14, iwr13 => iwr13, m13 => m13, m12 => m12, iwr12 => iwr12, clk4c => clk4c, iwr11 => iwr11, m11 => m11, m10 => m10, iwr10 => iwr10, iwr9 => iwr9, m9 => m9, m8 => m8, iwr8 => iwr8, iwr7 => iwr7, m7 => m7, m6 => m6, iwr6 => iwr6, iwr5 => iwr5, m5 => m5, m4 => m4, iwr4 => iwr4, iwr3 => iwr3, m3 => m3, m2 => m2, iwr2 => iwr2, iwr1 => iwr1, m1 => m1, m0 => m0, iwr0 => iwr0, iwr31 => iwr31, m31 => m31, m30 => m30, iwr30 => iwr30, iwr29 => iwr29, m29 => m29, m28 => m28, iwr28 => iwr28, iwr27 => iwr27, m27 => m27, m26 => m26, iwr26 => iwr26, iwr25 => iwr25, m25 => m25, m24 => m24, iwr24 => iwr24, iwr23 => iwr23, m23 => m23, m22 => m22, iwr22 => iwr22, iwr21 => iwr21, m21 => m21, m20 => m20, iwr20 => iwr20, iwr19 => iwr19, m19 => m19, m18 => m18, iwr18 => iwr18, iwr17 => iwr17, m17 => m17, m16 => m16, iwr16 => iwr16);
  i_pctl : entity icmem_book.pctl(ttl) port map(\-promenable\ => \-promenable\, gnd => gnd, i46 => i46, hi2 => hi2, pc0 => pc0, \-prompc0\ => \-prompc0\, pc1 => pc1, \-prompc1\ => \-prompc1\, pc2 => pc2, \-prompc2\ => \-prompc2\, \-prompc3\ => \-prompc3\, pc3 => pc3, \-prompc4\ => \-prompc4\, pc4 => pc4, pc9 => pc9, \-promce0\ => \-promce0\, \-prompc9\ => \-prompc9\, \-promce1\ => \-promce1\, \bottom.1k\ => \bottom.1k\, \-idebug\ => \-idebug\, \-promdisabled\ => \-promdisabled\, \-iwriteda\ => \-iwriteda\, pc13 => pc13, pc12 => pc12, pc11 => pc11, pc10 => pc10, pc5 => pc5, \-prompc5\ => \-prompc5\, pc6 => pc6, \-prompc6\ => \-prompc6\, pc7 => pc7, \-prompc7\ => \-prompc7\, \-prompc8\ => \-prompc8\, pc8 => pc8, \-ape\ => \-ape\, \-pdlpe\ => \-pdlpe\, \-spe\ => \-spe\, \-mpe\ => \-mpe\, tilt1 => tilt1, tilt0 => tilt0, \-mempe\ => \-mempe\, \-v1pe\ => \-v1pe\, \-v0pe\ => \-v0pe\, promenable => promenable, dpe => dpe, \-dpe\ => \-dpe\, ipe => ipe, \-ipe\ => \-ipe\);
  i_prom0 : entity icmem_book.prom0(ttl) port map(\-prompc0\ => \-prompc0\, \-prompc1\ => \-prompc1\, \-prompc2\ => \-prompc2\, \-prompc3\ => \-prompc3\, \-prompc4\ => \-prompc4\, i32 => i32, i33 => i33, i34 => i34, i35 => i35, i36 => i36, i37 => i37, i38 => i38, i39 => i39, \-promce0\ => \-promce0\, \-prompc5\ => \-prompc5\, \-prompc6\ => \-prompc6\, \-prompc7\ => \-prompc7\, \-prompc8\ => \-prompc8\, i40 => i40, i41 => i41, i42 => i42, i43 => i43, i44 => i44, i45 => i45, i47 => i47, i48 => i48, i24 => i24, i25 => i25, i26 => i26, i27 => i27, i28 => i28, i29 => i29, i30 => i30, i31 => i31, i16 => i16, i17 => i17, i18 => i18, i19 => i19, i20 => i20, i21 => i21, i22 => i22, i23 => i23, i0 => i0, i1 => i1, i2 => i2, i3 => i3, i4 => i4, i5 => i5, i6 => i6, i7 => i7, i8 => i8, i9 => i9, i10 => i10, i11 => i11, i12 => i12, i13 => i13, i14 => i14, i15 => i15);
  i_prom1 : entity icmem_book.prom1(ttl) port map(\-prompc0\ => \-prompc0\, \-prompc1\ => \-prompc1\, \-prompc2\ => \-prompc2\, \-prompc3\ => \-prompc3\, \-prompc4\ => \-prompc4\, i24 => i24, i25 => i25, i26 => i26, i27 => i27, i28 => i28, i29 => i29, i30 => i30, i31 => i31, \-promce1\ => \-promce1\, \-prompc5\ => \-prompc5\, \-prompc6\ => \-prompc6\, \-prompc7\ => \-prompc7\, \-prompc8\ => \-prompc8\, i32 => i32, i33 => i33, i34 => i34, i35 => i35, i36 => i36, i37 => i37, i38 => i38, i39 => i39, i40 => i40, i41 => i41, i42 => i42, i43 => i43, i44 => i44, i45 => i45, i47 => i47, i48 => i48, i16 => i16, i17 => i17, i18 => i18, i19 => i19, i20 => i20, i21 => i21, i22 => i22, i23 => i23, i0 => i0, i1 => i1, i2 => i2, i3 => i3, i4 => i4, i5 => i5, i6 => i6, i7 => i7, i8 => i8, i9 => i9, i10 => i10, i11 => i11, i12 => i12, i13 => i13, i14 => i14, i15 => i15);
  i_debug : entity icmem_book.debug(ttl) port map(\-idebug\ => \-idebug\, i39 => i39, spy7 => spy7, spy6 => spy6, i38 => i38, i37 => i37, spy5 => spy5, spy4 => spy4, i36 => i36, \-lddbirh\ => \-lddbirh\, i35 => i35, spy3 => spy3, spy2 => spy2, i34 => i34, i33 => i33, spy1 => spy1, spy0 => spy0, i32 => i32, i31 => i31, spy15 => spy15, spy14 => spy14, i30 => i30, i29 => i29, spy13 => spy13, spy12 => spy12, i28 => i28, \-lddbirm\ => \-lddbirm\, i27 => i27, spy11 => spy11, spy10 => spy10, i26 => i26, i25 => i25, spy9 => spy9, spy8 => spy8, i24 => i24, i23 => i23, i22 => i22, i21 => i21, i20 => i20, i19 => i19, i18 => i18, i17 => i17, i16 => i16, i15 => i15, i14 => i14, i13 => i13, i12 => i12, \-lddbirl\ => \-lddbirl\, i11 => i11, i10 => i10, i9 => i9, i8 => i8, i7 => i7, i6 => i6, i5 => i5, i4 => i4, i3 => i3, i2 => i2, i1 => i1, i0 => i0, i47 => i47, i46 => i46, i45 => i45, i44 => i44, i43 => i43, i42 => i42, i41 => i41, i40 => i40);


--- Microinstrction Modification and Main Instruction Register (ior)
  i_ior : entity cadr_book.ior(ttl) port map(i12 => i12, ob12 => ob12, iob12 => iob12, i13 => i13, ob13 => ob13, iob13 => iob13, iob14 => iob14, i14 => i14, ob14 => ob14, iob15 => iob15, i15 => i15, ob15 => ob15, i8 => i8, ob8 => ob8, iob8 => iob8, i9 => i9, ob9 => ob9, iob9 => iob9, iob10 => iob10, i10 => i10, ob10 => ob10, iob11 => iob11, i11 => i11, ob11 => ob11, i4 => i4, ob4 => ob4, iob4 => iob4, i5 => i5, ob5 => ob5, iob5 => iob5, iob6 => iob6, i6 => i6, ob6 => ob6, iob7 => iob7, i7 => i7, ob7 => ob7, i0 => i0, ob0 => ob0, iob0 => iob0, i1 => i1, ob1 => ob1, iob1 => iob1, iob2 => iob2, i2 => i2, ob2 => ob2, iob3 => iob3, i3 => i3, ob3 => ob3, i20 => i20, ob20 => ob20, iob20 => iob20, i21 => i21, ob21 => ob21, iob21 => iob21, iob22 => iob22, i22 => i22, ob22 => ob22, iob23 => iob23, i23 => i23, ob23 => ob23, i16 => i16, ob16 => ob16, iob16 => iob16, i17 => i17, ob17 => ob17, iob17 => iob17, iob18 => iob18, i18 => i18, ob18 => ob18, iob19 => iob19, i19 => i19, ob19 => ob19, i44 => i44, iob44 => iob44, i45 => i45, iob45 => iob45, iob46 => iob46, i46 => i46, iob47 => iob47, i47 => i47, i40 => i40, iob40 => iob40, i41 => i41, iob41 => iob41, iob42 => iob42, i42 => i42, iob43 => iob43, i43 => i43, i36 => i36, iob36 => iob36, i37 => i37, iob37 => iob37, iob38 => iob38, i38 => i38, iob39 => iob39, i39 => i39, i32 => i32, iob32 => iob32, i33 => i33, iob33 => iob33, iob34 => iob34, i34 => i34, iob35 => iob35, i35 => i35, i28 => i28, iob28 => iob28, i29 => i29, iob29 => iob29, iob30 => iob30, i30 => i30, iob31 => iob31, i31 => i31, i24 => i24, ob24 => ob24, iob24 => iob24, i25 => i25, ob25 => ob25, iob25 => iob25, iob26 => iob26, i26 => i26, iob27 => iob27, i27 => i27);
  i_ireg : entity cadr_book.ireg(ttl) port map(\-destimod0\ => \-destimod0\, ir15 => ir15, iob15 => iob15, i15 => i15, i14 => i14, iob14 => iob14, ir14 => ir14, clk3a => clk3a, ir13 => ir13, iob13 => iob13, i13 => i13, i12 => i12, iob12 => iob12, ir12 => ir12, ir11 => ir11, iob11 => iob11, i11 => i11, i10 => i10, iob10 => iob10, ir10 => ir10, ir9 => ir9, iob9 => iob9, i9 => i9, i8 => i8, iob8 => iob8, ir8 => ir8, ir7 => ir7, iob7 => iob7, i7 => i7, i6 => i6, iob6 => iob6, ir6 => ir6, ir5 => ir5, iob5 => iob5, i5 => i5, i4 => i4, iob4 => iob4, ir4 => ir4, ir3 => ir3, iob3 => iob3, i3 => i3, i2 => i2, iob2 => iob2, ir2 => ir2, ir1 => ir1, iob1 => iob1, i1 => i1, i0 => i0, iob0 => iob0, ir0 => ir0, ir23 => ir23, iob23 => iob23, i23 => i23, i22 => i22, iob22 => iob22, ir22 => ir22, clk3b => clk3b, ir21 => ir21, iob21 => iob21, i21 => i21, i20 => i20, iob20 => iob20, ir20 => ir20, ir19 => ir19, iob19 => iob19, i19 => i19, i18 => i18, iob18 => iob18, ir18 => ir18, ir17 => ir17, iob17 => iob17, i17 => i17, i16 => i16, iob16 => iob16, ir16 => ir16, \-destimod1\ => \-destimod1\, i48 => i48, gnd => gnd, ir48 => ir48, ir47 => ir47, iob47 => iob47, i47 => i47, i46 => i46, iob46 => iob46, ir46 => ir46, ir45 => ir45, iob45 => iob45, i45 => i45, i44 => i44, iob44 => iob44, ir44 => ir44, ir43 => ir43, iob43 => iob43, i43 => i43, i42 => i42, iob42 => iob42, ir42 => ir42, ir41 => ir41, iob41 => iob41, i41 => i41, i40 => i40, iob40 => iob40, ir40 => ir40, ir39 => ir39, iob39 => iob39, i39 => i39, i38 => i38, iob38 => iob38, ir38 => ir38, ir37 => ir37, iob37 => iob37, i37 => i37, i36 => i36, iob36 => iob36, ir36 => ir36, ir35 => ir35, iob35 => iob35, i35 => i35, i34 => i34, iob34 => iob34, ir34 => ir34, ir33 => ir33, iob33 => iob33, i33 => i33, i32 => i32, iob32 => iob32, ir32 => ir32, ir31 => ir31, iob31 => iob31, i31 => i31, i30 => i30, iob30 => iob30, ir30 => ir30, ir29 => ir29, iob29 => iob29, i29 => i29, i28 => i28, iob28 => iob28, ir28 => ir28, ir27 => ir27, iob27 => iob27, i27 => i27, i26 => i26, iob26 => iob26, ir26 => ir26, ir25 => ir25, iob25 => iob25, i25 => i25, i24 => i24, iob24 => iob24, ir24 => ir24);


--- IR Decoding (source?)
  i_source : entity cadr_book.source(ttl) port map(\-iralu\ => \-iralu\, \-irbyte\ => \-irbyte\, dest => dest, \-destmem\ => \-destmem\, ir23 => ir23, destm => destm, \-specalu\ => \-specalu\, ir8 => ir8, iralu => iralu, ir22 => ir22, \-ir22\ => \-ir22\, ir25 => ir25, \-ir25\ => \-ir25\, irdisp => irdisp, \-irdisp\ => \-irdisp\, irjump => irjump, \-irjump\ => \-irjump\, ir3 => ir3, ir4 => ir4, \-mul\ => \-mul\, \-div\ => \-div\, nop => nop, ir43 => ir43, ir44 => ir44, \-funct3\ => \-funct3\, \-funct2\ => \-funct2\, \-funct1\ => \-funct1\, \-funct0\ => \-funct0\, ir11 => ir11, ir10 => ir10, ir19 => ir19, ir20 => ir20, ir21 => ir21, \-destintctl\ => \-destintctl\, \-destlc\ => \-destlc\, \-destimod1\ => \-destimod1\, \-destimod0\ => \-destimod0\, \-destspc\ => \-destspc\, \-destpdlp\ => \-destpdlp\, \-destpdlx\ => \-destpdlx\, \-destpdl(x)\ => \-destpdl(x)\, \-destpdl(p)\ => \-destpdl(p)\, \-destpdltop\ => \-destpdltop\, ir26 => ir26, ir27 => ir27, ir28 => ir28, \-ir31\ => \-ir31\, ir29 => ir29, hi5 => hi5, \-srcq\ => \-srcq\, \-srcopc\ => \-srcopc\, \-srcpdltop\ => \-srcpdltop\, \-srcpdlpop\ => \-srcpdlpop\, \-srcpdlidx\ => \-srcpdlidx\, \-srcpdlptr\ => \-srcpdlptr\, \-srcspc\ => \-srcspc\, \-srcdc\ => \-srcdc\, gnd => gnd, \-srcspcpop\ => \-srcspcpop\, \-srclc\ => \-srclc\, \-srcmd\ => \-srcmd\, \-srcmap\ => \-srcmap\, \-srcvma\ => \-srcvma\, \destimod0_l\ => \destimod0_l\, \iwrited_l\ => \iwrited_l\, \-destmdr\ => \-destmdr\, \-destvma\ => \-destvma\, \-idebug\ => \-idebug\, imod => imod);


--- A Memory (amem)
  i_actl : entity cadr_book.actl(ttl) port map(clk3e => clk3e, wadr0 => wadr0, ir32 => ir32, \-aadr0b\ => \-aadr0b\, wadr1 => wadr1, ir33 => ir33, \-aadr1b\ => \-aadr1b\, \-aadr2b\ => \-aadr2b\, ir34 => ir34, wadr2 => wadr2, \-aadr3b\ => \-aadr3b\, ir35 => ir35, wadr3 => wadr3, gnd => gnd, clk3d => clk3d, wadr4 => wadr4, ir36 => ir36, \-aadr4b\ => \-aadr4b\, wadr5 => wadr5, ir37 => ir37, \-aadr5b\ => \-aadr5b\, \-aadr6b\ => \-aadr6b\, ir38 => ir38, wadr6 => wadr6, \-aadr7b\ => \-aadr7b\, ir39 => ir39, wadr7 => wadr7, \-aadr0a\ => \-aadr0a\, \-aadr1a\ => \-aadr1a\, \-aadr2a\ => \-aadr2a\, \-aadr3a\ => \-aadr3a\, \-aadr4a\ => \-aadr4a\, \-aadr5a\ => \-aadr5a\, \-aadr6a\ => \-aadr6a\, \-aadr7a\ => \-aadr7a\, wadr8 => wadr8, ir40 => ir40, \-aadr8a\ => \-aadr8a\, wadr9 => wadr9, ir41 => ir41, \-aadr9a\ => \-aadr9a\, \-aadr8b\ => \-aadr8b\, \-aadr9b\ => \-aadr9b\, apass1 => apass1, apass2 => apass2, \-apass\ => \-apass\, tse3a => tse3a, \-amemenb\ => \-amemenb\, hi3 => hi3, \-reset\ => \-reset\, ir14 => ir14, ir15 => ir15, ir16 => ir16, ir17 => ir17, destmd => destmd, destm => destm, dest => dest, destd => destd, ir21 => ir21, ir20 => ir20, ir19 => ir19, ir18 => ir18, ir23 => ir23, ir22 => ir22, wp3a => wp3a, \-awpa\ => \-awpa\, \-awpb\ => \-awpb\, \-awpc\ => \-awpc\, tse4a => tse4a, apassenb => apassenb, \-apassenb\ => \-apassenb\);
  i_amem0 : entity cadr_book.amem0(ttl) port map(gnd => gnd, \-aadr0b\ => \-aadr0b\, \-aadr1b\ => \-aadr1b\, \-aadr2b\ => \-aadr2b\, \-aadr3b\ => \-aadr3b\, \-aadr4b\ => \-aadr4b\, amem22 => amem22, \-aadr5b\ => \-aadr5b\, \-aadr6b\ => \-aadr6b\, \-aadr7b\ => \-aadr7b\, \-aadr8b\ => \-aadr8b\, \-aadr9b\ => \-aadr9b\, \-awpa\ => \-awpa\, l22 => l22, amem20 => amem20, l20 => l20, amem18 => amem18, l18 => l18, amem16 => amem16, l16 => l16, amem23 => amem23, l23 => l23, amem21 => amem21, l21 => l21, amem19 => amem19, l19 => l19, amem17 => amem17, l17 => l17, amemparity => amemparity, lparity => lparity, amem30 => amem30, l30 => l30, amem28 => amem28, l28 => l28, amem26 => amem26, l26 => l26, amem24 => amem24, l24 => l24, amem31 => amem31, l31 => l31, amem29 => amem29, l29 => l29, amem27 => amem27, l27 => l27, amem25 => amem25, l25 => l25);
  i_amem1 : entity cadr_book.amem1(ttl) port map(gnd => gnd, \-aadr0a\ => \-aadr0a\, \-aadr1a\ => \-aadr1a\, \-aadr2a\ => \-aadr2a\, \-aadr3a\ => \-aadr3a\, \-aadr4a\ => \-aadr4a\, amem6 => amem6, \-aadr5a\ => \-aadr5a\, \-aadr6a\ => \-aadr6a\, \-aadr7a\ => \-aadr7a\, \-aadr8a\ => \-aadr8a\, \-aadr9a\ => \-aadr9a\, \-awpc\ => \-awpc\, l6 => l6, amem4 => amem4, l4 => l4, amem2 => amem2, l2 => l2, amem0 => amem0, l0 => l0, amem7 => amem7, l7 => l7, amem5 => amem5, l5 => l5, amem3 => amem3, l3 => l3, amem1 => amem1, l1 => l1, amem14 => amem14, \-awpb\ => \-awpb\, l14 => l14, amem12 => amem12, l12 => l12, amem10 => amem10, l10 => l10, amem8 => amem8, l8 => l8, amem15 => amem15, l15 => l15, amem13 => amem13, l13 => l13, amem11 => amem11, l11 => l11, amem9 => amem9, l9 => l9);
  i_alatch : entity cadr_book.alatch(ttl) port map(\-amemenb\ => \-amemenb\, a23 => a23, amem23 => amem23, amem22 => amem22, a22 => a22, a21 => a21, amem21 => amem21, amem20 => amem20, a20 => a20, clk3e => clk3e, a19 => a19, amem19 => amem19, amem18 => amem18, a18 => a18, a17 => a17, amem17 => amem17, amem16 => amem16, a16 => a16, \-apassenb\ => \-apassenb\, l15 => l15, a8 => a8, l14 => l14, a9 => a9, l13 => l13, a10 => a10, l12 => l12, a11 => a11, l11 => l11, a12 => a12, l10 => l10, a13 => a13, l9 => l9, a14 => a14, l8 => l8, a15 => a15, apassenb => apassenb, amem15 => amem15, amem14 => amem14, amem13 => amem13, amem12 => amem12, amem11 => amem11, amem10 => amem10, amem9 => amem9, amem8 => amem8, l7 => l7, a0 => a0, l6 => l6, a1 => a1, l5 => l5, a2 => a2, l4 => l4, a3 => a3, l3 => l3, a4 => a4, l2 => l2, a5 => a5, l1 => l1, a6 => a6, l0 => l0, a7 => a7, amem7 => amem7, amem6 => amem6, amem5 => amem5, amem4 => amem4, amem3 => amem3, amem2 => amem2, amem1 => amem1, amem0 => amem0, hi5 => hi5, a31b => a31b, aparity => aparity, lparity => lparity, l31 => l31, amemparity => amemparity, amem31 => amem31, a24 => a24, l30 => l30, a25 => a25, l29 => l29, a26 => a26, l28 => l28, a27 => a27, l27 => l27, a28 => a28, l26 => l26, a29 => a29, l25 => l25, a30 => a30, l24 => l24, a31a => a31a, amem30 => amem30, amem29 => amem29, amem28 => amem28, amem27 => amem27, amem26 => amem26, amem25 => amem25, amem24 => amem24, l23 => l23, l22 => l22, l21 => l21, l20 => l20, l19 => l19, l18 => l18, l17 => l17, l16 => l16);
  i_apar : entity cadr_book.apar(ttl) port map(a26 => a26, a27 => a27, a28 => a28, a29 => a29, a30 => a30, a31b => a31b, aparity => aparity, aparok => aparok, aparl => aparl, aparm => aparm, gnd => gnd, a24 => a24, a25 => a25, a17 => a17, a18 => a18, a19 => a19, a20 => a20, a21 => a21, a22 => a22, a23 => a23, a12 => a12, a13 => a13, a14 => a14, a15 => a15, a16 => a16, a5 => a5, a6 => a6, a7 => a7, a8 => a8, a9 => a9, a10 => a10, a11 => a11, a0 => a0, a1 => a1, a2 => a2, a3 => a3, a4 => a4, m17 => m17, m18 => m18, m19 => m19, m20 => m20, m21 => m21, m22 => m22, m23 => m23, mparm => mparm, m12 => m12, m13 => m13, m14 => m14, m15 => m15, m16 => m16, m5 => m5, m6 => m6, m7 => m7, m8 => m8, m9 => m9, m10 => m10, m11 => m11, mparl => mparl, m0 => m0, m1 => m1, m2 => m2, m3 => m3, m4 => m4, mpareven => mpareven, srcm => srcm, mmemparok => mmemparok, pdlenb => pdlenb, pdlparok => pdlparok, m26 => m26, m27 => m27, m28 => m28, m29 => m29, m30 => m30, m31 => m31, mparity => mparity, mparodd => mparodd, m24 => m24, m25 => m25);


--- M Memory (mmem)
  i_mctl : entity cadr_book.mctl(ttl) port map(clk4e => clk4e, wadr4 => wadr4, ir30 => ir30, \-madr4a\ => \-madr4a\, \-madr4b\ => \-madr4b\, gnd => gnd, wadr0 => wadr0, ir26 => ir26, \-madr0b\ => \-madr0b\, wadr1 => wadr1, ir27 => ir27, \-madr1b\ => \-madr1b\, \-madr2b\ => \-madr2b\, ir28 => ir28, wadr2 => wadr2, \-madr3b\ => \-madr3b\, ir29 => ir29, wadr3 => wadr3, mmem15 => mmem15, mmem14 => mmem14, mmem13 => mmem13, mmem12 => mmem12, mmem11 => mmem11, mmem10 => mmem10, mmem9 => mmem9, mmem8 => mmem8, mmem7 => mmem7, mmem6 => mmem6, mmem5 => mmem5, mmem4 => mmem4, mmem3 => mmem3, mmem2 => mmem2, mmem1 => mmem1, mmem0 => mmem0, mpass => mpass, tse4a => tse4a, srcm => srcm, hi2 => hi2, \-ir31\ => \-ir31\, \-mpass\ => \-mpass\, mpassl => mpassl, \-mpassm\ => \-mpassm\, \-mpassl\ => \-mpassl\, destmd => destmd, \-madr0a\ => \-madr0a\, \-madr1a\ => \-madr1a\, \-madr2a\ => \-madr2a\, \-madr3a\ => \-madr3a\, mmemparity => mmemparity, mmem31 => mmem31, mmem30 => mmem30, mmem29 => mmem29, mmem28 => mmem28, mmem27 => mmem27, mmem26 => mmem26, mmem25 => mmem25, mmem24 => mmem24, mmem23 => mmem23, mmem22 => mmem22, mmem21 => mmem21, mmem20 => mmem20, mmem19 => mmem19, mmem18 => mmem18, mmem17 => mmem17, mmem16 => mmem16, wp4b => wp4b, \-mwpa\ => \-mwpa\, \-mwpb\ => \-mwpb\);
  i_mmem : entity cadr_book.mmem(ttl) port map(\-mwpa\ => \-mwpa\, gnd => gnd, l16 => l16, \-madr4a\ => \-madr4a\, hi3 => hi3, mmem16 => mmem16, mmem17 => mmem17, \-madr3a\ => \-madr3a\, \-madr2a\ => \-madr2a\, \-madr1a\ => \-madr1a\, \-madr0a\ => \-madr0a\, l17 => l17, \-mwpb\ => \-mwpb\, l12 => l12, \-madr4b\ => \-madr4b\, hi2 => hi2, mmem12 => mmem12, mmem13 => mmem13, \-madr3b\ => \-madr3b\, \-madr2b\ => \-madr2b\, \-madr1b\ => \-madr1b\, \-madr0b\ => \-madr0b\, l13 => l13, l8 => l8, mmem8 => mmem8, mmem9 => mmem9, l9 => l9, l4 => l4, mmem4 => mmem4, mmem5 => mmem5, l5 => l5, l0 => l0, mmem0 => mmem0, mmem1 => mmem1, l1 => l1, l18 => l18, mmem18 => mmem18, mmem19 => mmem19, l19 => l19, l14 => l14, mmem14 => mmem14, mmem15 => mmem15, l15 => l15, l10 => l10, mmem10 => mmem10, mmem11 => mmem11, l11 => l11, l6 => l6, mmem6 => mmem6, mmem7 => mmem7, l7 => l7, l2 => l2, mmem2 => mmem2, mmem3 => mmem3, l3 => l3, l28 => l28, mmem28 => mmem28, mmem29 => mmem29, l29 => l29, l24 => l24, mmem24 => mmem24, mmem25 => mmem25, l25 => l25, l20 => l20, mmem20 => mmem20, mmem21 => mmem21, l21 => l21, lparity => lparity, mmemparity => mmemparity, l30 => l30, mmem30 => mmem30, mmem31 => mmem31, l31 => l31, l26 => l26, mmem26 => mmem26, mmem27 => mmem27, l27 => l27, l22 => l22, mmem22 => mmem22, mmem23 => mmem23, l23 => l23);
  i_mlatch : entity cadr_book.mlatch(ttl) port map(\-mpassm\ => \-mpassm\, m23 => m23, mmem23 => mmem23, mmem22 => mmem22, m22 => m22, m21 => m21, mmem21 => mmem21, mmem20 => mmem20, m20 => m20, clk4a => clk4a, m19 => m19, mmem19 => mmem19, mmem18 => mmem18, m18 => m18, m17 => m17, mmem17 => mmem17, mmem16 => mmem16, m16 => m16, m15 => m15, mmem15 => mmem15, mmem14 => mmem14, m14 => m14, m13 => m13, mmem13 => mmem13, mmem12 => mmem12, m12 => m12, m11 => m11, mmem11 => mmem11, mmem10 => mmem10, m10 => m10, m9 => m9, mmem9 => mmem9, mmem8 => mmem8, m8 => m8, m7 => m7, mmem7 => mmem7, mmem6 => mmem6, m6 => m6, m5 => m5, mmem5 => mmem5, mmem4 => mmem4, m4 => m4, m3 => m3, mmem3 => mmem3, mmem2 => mmem2, m2 => m2, m1 => m1, mmem1 => mmem1, mmem0 => mmem0, m0 => m0, \-mpassl\ => \-mpassl\, l15 => l15, mf8 => mf8, l14 => l14, mf9 => mf9, l13 => l13, mf10 => mf10, l12 => l12, mf11 => mf11, l11 => l11, mf12 => mf12, l10 => l10, mf13 => mf13, l9 => l9, mf14 => mf14, l8 => l8, mf15 => mf15, mpassl => mpassl, l7 => l7, mf0 => mf0, l6 => l6, mf1 => mf1, l5 => l5, mf2 => mf2, l4 => l4, mf3 => mf3, l3 => l3, mf4 => mf4, l2 => l2, mf5 => mf5, l1 => l1, mf6 => mf6, l0 => l0, mf7 => mf7, mmemparity => mmemparity, mparity => mparity, m31 => m31, mmem31 => mmem31, mmem30 => mmem30, m30 => m30, m29 => m29, mmem29 => mmem29, mmem28 => mmem28, m28 => m28, m27 => m27, mmem27 => mmem27, mmem26 => mmem26, m26 => m26, m25 => m25, mmem25 => mmem25, mmem24 => mmem24, m24 => m24, l31 => l31, mf24 => mf24, l30 => l30, mf25 => mf25, l29 => l29, mf26 => mf26, l28 => l28, mf27 => mf27, l27 => l27, mf28 => mf28, l26 => l26, mf29 => mf29, l25 => l25, mf30 => mf30, l24 => l24, mf31 => mf31, l23 => l23, mf16 => mf16, l22 => l22, mf17 => mf17, l21 => l21, mf18 => mf18, l20 => l20, mf19 => mf19, l19 => l19, mf20 => mf20, l18 => l18, mf21 => mf21, l17 => l17, mf22 => mf22, l16 => l16, mf23 => mf23);
  i_mf : entity cadr_book.mf(ttl) port map(tse1a => tse1a, mfenb => mfenb, \-mfdrive\ => \-mfdrive\, mf23 => mf23, m16 => m16, mf22 => mf22, m17 => m17, mf21 => mf21, m18 => m18, mf20 => mf20, m19 => m19, mf19 => mf19, m20 => m20, mf18 => mf18, m21 => m21, mf17 => mf17, m22 => m22, mf16 => mf16, m23 => m23, mfdrive => mfdrive, mf15 => mf15, m8 => m8, mf14 => mf14, m9 => m9, mf13 => mf13, m10 => m10, mf12 => mf12, m11 => m11, mf11 => mf11, m12 => m12, mf10 => mf10, m13 => m13, mf9 => mf9, m14 => m14, mf8 => mf8, m15 => m15, mf7 => mf7, m0 => m0, mf6 => mf6, m1 => m1, mf5 => mf5, m2 => m2, mf4 => mf4, m3 => m3, mf3 => mf3, m4 => m4, mf2 => mf2, m5 => m5, mf1 => mf1, m6 => m6, mf0 => mf0, m7 => m7, mf31 => mf31, m24 => m24, mf30 => mf30, m25 => m25, mf29 => mf29, m26 => m26, mf28 => mf28, m27 => m27, mf27 => mf27, m28 => m28, mf26 => mf26, m29 => m29, mf25 => mf25, m30 => m30, mf24 => mf24, m31 => m31, pdlenb => pdlenb, spcenb => spcenb, \-srcm\ => \-srcm\, \-ir31\ => \-ir31\, \-mpass\ => \-mpass\);


--- Stack Buffer (pdl)
  i_pdlptr : entity cadr_book.pdlptr(ttl) port map(\-srcpdlpop\ => \-srcpdlpop\, clk3f => clk3f, ob8 => ob8, ob9 => ob9, gnd => gnd, \-destpdlp\ => \-destpdlp\, \-pdlcry7\ => \-pdlcry7\, pdlptr9 => pdlptr9, pdlptr8 => pdlptr8, \-destpdlx\ => \-destpdlx\, pdlidx6 => pdlidx6, ob6 => ob6, ob7 => ob7, pdlidx7 => pdlidx7, pdlidx8 => pdlidx8, pdlidx9 => pdlidx9, ob4 => ob4, ob5 => ob5, \-pdlcry3\ => \-pdlcry3\, pdlptr7 => pdlptr7, pdlptr6 => pdlptr6, pdlptr5 => pdlptr5, pdlptr4 => pdlptr4, pdlidx0 => pdlidx0, ob0 => ob0, ob1 => ob1, pdlidx1 => pdlidx1, ob2 => ob2, pdlidx2 => pdlidx2, pdlidx3 => pdlidx3, ob3 => ob3, pdlidx4 => pdlidx4, pdlidx5 => pdlidx5, \-pdlcnt\ => \-pdlcnt\, pdlptr3 => pdlptr3, pdlptr2 => pdlptr2, pdlptr1 => pdlptr1, pdlptr0 => pdlptr0, \-ppdrive\ => \-ppdrive\, mf0 => mf0, mf1 => mf1, mf2 => mf2, mf3 => mf3, pidrive => pidrive, mf8 => mf8, mf9 => mf9, mf10 => mf10, mf11 => mf11, mf4 => mf4, mf5 => mf5, mf6 => mf6, mf7 => mf7, srcpdlidx => srcpdlidx, tse4b => tse4b, srcpdlptr => srcpdlptr);
  i_pdlctl : entity cadr_book.pdlctl(ttl) port map(\-reset\ => \-reset\, pdlwrited => pdlwrited, \-pdlwrited\ => \-pdlwrited\, pdlwrite => pdlwrite, \-destpdl(x)\ => \-destpdl(x)\, pwidx => pwidx, \-pwidx\ => \-pwidx\, clk4f => clk4f, imodd => imodd, \-imodd\ => \-imodd\, imod => imod, \-destspc\ => \-destspc\, \-destspcd\ => \-destspcd\, \-pdlpb\ => \-pdlpb\, pdlptr0 => pdlptr0, pdlidx0 => pdlidx0, \-pdla0b\ => \-pdla0b\, pdlptr1 => pdlptr1, pdlidx1 => pdlidx1, \-pdla1b\ => \-pdla1b\, \-pdla2b\ => \-pdla2b\, pdlidx2 => pdlidx2, pdlptr2 => pdlptr2, \-pdla3b\ => \-pdla3b\, pdlidx3 => pdlidx3, pdlptr3 => pdlptr3, gnd => gnd, \-pdlpa\ => \-pdlpa\, pdlptr8 => pdlptr8, pdlidx8 => pdlidx8, \-pdla8b\ => \-pdla8b\, pdlptr9 => pdlptr9, pdlidx9 => pdlidx9, \-pdla9b\ => \-pdla9b\, \-pdla0a\ => \-pdla0a\, \-pdla1a\ => \-pdla1a\, \-pdla2a\ => \-pdla2a\, \-pdla3a\ => \-pdla3a\, \-pdla4a\ => \-pdla4a\, pdlidx4 => pdlidx4, pdlptr4 => pdlptr4, \-pdla5a\ => \-pdla5a\, pdlidx5 => pdlidx5, pdlptr5 => pdlptr5, \-destpdl(p)\ => \-destpdl(p)\, \-pdlcnt\ => \-pdlcnt\, clk4b => clk4b, ir30 => ir30, \-clk4e\ => \-clk4e\, \-srcpdlpop\ => \-srcpdlpop\, \-srcpdltop\ => \-srcpdltop\, pdlenb => pdlenb, tse4b => tse4b, \-pdldrive\ => \-pdldrive\, \-destpdltop\ => \-destpdltop\, \-pdla4b\ => \-pdla4b\, \-pdla5b\ => \-pdla5b\, \-pdla6b\ => \-pdla6b\, pdlidx6 => pdlidx6, pdlptr6 => pdlptr6, \-pdla7b\ => \-pdla7b\, pdlidx7 => pdlidx7, pdlptr7 => pdlptr7, wp4a => wp4a, \-pwpa\ => \-pwpa\, \-pwpb\ => \-pwpb\, \-pwpc\ => \-pwpc\, \-pdla6a\ => \-pdla6a\, \-pdla7a\ => \-pdla7a\, \-pdla8a\ => \-pdla8a\, \-pdla9a\ => \-pdla9a\, nop => nop);
  i_pdl0 : entity cadr_book.pdl0(ttl) port map(gnd => gnd, \-pdla0b\ => \-pdla0b\, \-pdla1b\ => \-pdla1b\, \-pdla2b\ => \-pdla2b\, \-pdla3b\ => \-pdla3b\, \-pdla4b\ => \-pdla4b\, pdlparity => pdlparity, \-pdla5b\ => \-pdla5b\, \-pdla6b\ => \-pdla6b\, \-pdla7b\ => \-pdla7b\, \-pdla8b\ => \-pdla8b\, \-pdla9b\ => \-pdla9b\, \-pwpa\ => \-pwpa\, lparity => lparity, pdl28 => pdl28, l28 => l28, pdl27 => pdl27, l27 => l27, pdl26 => pdl26, l26 => l26, pdl21 => pdl21, \-pwpb\ => \-pwpb\, l21 => l21, pdl20 => pdl20, l20 => l20, pdl19 => pdl19, l19 => l19, pdl18 => pdl18, l18 => l18, pdl31 => pdl31, l31 => l31, pdl30 => pdl30, l30 => l30, pdl29 => pdl29, l29 => l29, pdl25 => pdl25, l25 => l25, pdl24 => pdl24, l24 => l24, pdl23 => pdl23, l23 => l23, pdl22 => pdl22, l22 => l22, pdl17 => pdl17, l17 => l17, pdl16 => pdl16, l16 => l16);
  i_pdl1 : entity cadr_book.pdl1(ttl) port map(gnd => gnd, \-pdla0a\ => \-pdla0a\, \-pdla1a\ => \-pdla1a\, \-pdla2a\ => \-pdla2a\, \-pdla3a\ => \-pdla3a\, \-pdla4a\ => \-pdla4a\, pdl13 => pdl13, \-pdla5a\ => \-pdla5a\, \-pdla6a\ => \-pdla6a\, \-pdla7a\ => \-pdla7a\, \-pdla8a\ => \-pdla8a\, \-pdla9a\ => \-pdla9a\, \-pwpb\ => \-pwpb\, l13 => l13, pdl12 => pdl12, l12 => l12, pdl11 => pdl11, l11 => l11, pdl10 => pdl10, \-pwpc\ => \-pwpc\, l10 => l10, pdl4 => pdl4, l4 => l4, pdl3 => pdl3, l3 => l3, pdl2 => pdl2, l2 => l2, pdl1 => pdl1, l1 => l1, pdl0 => pdl0, l0 => l0, pdl15 => pdl15, l15 => l15, pdl14 => pdl14, l14 => l14, pdl9 => pdl9, l9 => l9, pdl8 => pdl8, l8 => l8, pdl7 => pdl7, l7 => l7, pdl6 => pdl6, l6 => l6, pdl5 => pdl5, l5 => l5);
  i_platch : entity cadr_book.platch(ttl) port map(\-pdldrive\ => \-pdldrive\, m15 => m15, pdl15 => pdl15, pdl14 => pdl14, m14 => m14, m13 => m13, pdl13 => pdl13, pdl12 => pdl12, m12 => m12, clk4a => clk4a, m11 => m11, pdl11 => pdl11, pdl10 => pdl10, m10 => m10, m9 => m9, pdl9 => pdl9, pdl8 => pdl8, m8 => m8, m7 => m7, pdl7 => pdl7, pdl6 => pdl6, m6 => m6, m5 => m5, pdl5 => pdl5, pdl4 => pdl4, m4 => m4, m3 => m3, pdl3 => pdl3, pdl2 => pdl2, m2 => m2, m1 => m1, pdl1 => pdl1, pdl0 => pdl0, m0 => m0, m31 => m31, pdl31 => pdl31, pdl30 => pdl30, m30 => m30, m29 => m29, pdl29 => pdl29, pdl28 => pdl28, m28 => m28, m27 => m27, pdl27 => pdl27, pdl26 => pdl26, m26 => m26, m25 => m25, pdl25 => pdl25, pdl24 => pdl24, m24 => m24, m23 => m23, pdl23 => pdl23, pdl22 => pdl22, m22 => m22, m21 => m21, pdl21 => pdl21, pdl20 => pdl20, m20 => m20, m19 => m19, pdl19 => pdl19, pdl18 => pdl18, m18 => m18, m17 => m17, pdl17 => pdl17, pdl16 => pdl16, m16 => m16, pdlparity => pdlparity, mparity => mparity);


--- The Shifter\Masker (sm)
  i_smctl : entity cadr_book.smctl(ttl) port map(\-sh4\ => \-sh4\, \-sr\ => \-sr\, \-s4\ => \-s4\, \-mr\ => \-mr\, \-irbyte\ => \-irbyte\, ir13 => ir13, ir12 => ir12, \-ir0\ => \-ir0\, s0 => s0, \-ir1\ => \-ir1\, s1 => s1, mskl4 => mskl4, ir9 => ir9, mskr4 => mskr4, mskl3cry => mskl3cry, s3a => s3a, \-sh3\ => \-sh3\, s3b => s3b, \-ir2\ => \-ir2\, s2a => s2a, s2b => s2b, s4 => s4, mskr0 => mskr0, mskr1 => mskr1, mskr2 => mskr2, mskl1 => mskl1, ir6 => ir6, mskl0 => mskl0, ir5 => ir5, gnd => gnd, mskl3 => mskl3, mskr3 => mskr3, ir8 => ir8, mskl2 => mskl2, ir7 => ir7);
  i_shift0 : entity cadr_book.shift0(ttl) port map(m5 => m5, m6 => m6, m7 => m7, m8 => m8, m9 => m9, m10 => m10, m11 => m11, s1 => s1, s0 => s0, sa11 => sa11, sa10 => sa10, gnd => gnd, sa9 => sa9, sa8 => sa8, m29 => m29, m30 => m30, m31 => m31, m0 => m0, m1 => m1, m2 => m2, m3 => m3, sa3 => sa3, sa2 => sa2, sa1 => sa1, sa0 => sa0, m12 => m12, m13 => m13, m14 => m14, m15 => m15, sa15 => sa15, sa14 => sa14, sa13 => sa13, sa12 => sa12, m4 => m4, sa7 => sa7, sa6 => sa6, sa5 => sa5, sa4 => sa4, sa18 => sa18, sa22 => sa22, sa26 => sa26, sa30 => sa30, s3a => s3a, s2a => s2a, r14 => r14, r10 => r10, \-s4\ => \-s4\, r6 => r6, r2 => r2, s4 => s4, sa19 => sa19, sa23 => sa23, sa27 => sa27, sa31 => sa31, r15 => r15, r11 => r11, r7 => r7, r3 => r3, sa16 => sa16, sa20 => sa20, sa24 => sa24, sa28 => sa28, r12 => r12, r8 => r8, r4 => r4, r0 => r0, sa17 => sa17, sa21 => sa21, sa25 => sa25, sa29 => sa29, r13 => r13, r9 => r9, r5 => r5, r1 => r1);
  i_shift1 : entity cadr_book.shift1(ttl) port map(m21 => m21, m22 => m22, m23 => m23, m24 => m24, m25 => m25, m26 => m26, m27 => m27, s1 => s1, s0 => s0, sa27 => sa27, sa26 => sa26, gnd => gnd, sa25 => sa25, sa24 => sa24, m13 => m13, m14 => m14, m15 => m15, m16 => m16, m17 => m17, m18 => m18, m19 => m19, sa19 => sa19, sa18 => sa18, sa17 => sa17, sa16 => sa16, m28 => m28, m29 => m29, m30 => m30, m31 => m31, sa31 => sa31, sa30 => sa30, sa29 => sa29, sa28 => sa28, m20 => m20, sa23 => sa23, sa22 => sa22, sa21 => sa21, sa20 => sa20, sa2 => sa2, sa6 => sa6, sa10 => sa10, sa14 => sa14, s3b => s3b, s2b => s2b, r30 => r30, r26 => r26, \-s4\ => \-s4\, r22 => r22, r18 => r18, s4 => s4, sa3 => sa3, sa7 => sa7, sa11 => sa11, sa15 => sa15, r31 => r31, r27 => r27, r23 => r23, r19 => r19, sa0 => sa0, sa4 => sa4, sa8 => sa8, sa12 => sa12, r28 => r28, r24 => r24, r20 => r20, r16 => r16, sa1 => sa1, sa5 => sa5, sa9 => sa9, sa13 => sa13, r29 => r29, r25 => r25, r21 => r21, r17 => r17);
  i_mskg4 : entity cadr_book.mskg4(ttl) port map(msk24 => msk24, msk25 => msk25, msk26 => msk26, msk27 => msk27, msk28 => msk28, msk29 => msk29, msk30 => msk30, msk31 => msk31, mskl0 => mskl0, mskl1 => mskl1, mskl2 => mskl2, mskl3 => mskl3, mskl4 => mskl4, gnd => gnd, mskr0 => mskr0, mskr1 => mskr1, mskr2 => mskr2, mskr3 => mskr3, mskr4 => mskr4, msk8 => msk8, msk9 => msk9, msk10 => msk10, msk11 => msk11, msk12 => msk12, msk13 => msk13, msk14 => msk14, msk15 => msk15, ir31 => ir31, \-ir31\ => \-ir31\, ir13 => ir13, \-ir13\ => \-ir13\, \-ir12\ => \-ir12\, ir12 => ir12, msk16 => msk16, msk17 => msk17, msk18 => msk18, msk19 => msk19, msk20 => msk20, msk21 => msk21, msk22 => msk22, msk23 => msk23, aeqm => aeqm, msk0 => msk0, msk1 => msk1, msk2 => msk2, msk3 => msk3, msk4 => msk4, msk5 => msk5, msk6 => msk6, msk7 => msk7);


--- The ALU (alu)
  i_aluc4 : entity cadr_book.aluc4(ttl) port map(\-aluf0\ => \-aluf0\, aluf0b => aluf0b, \-aluf1\ => \-aluf1\, aluf1b => aluf1b, aluf2b => aluf2b, \-aluf2\ => \-aluf2\, aluf3b => aluf3b, \-aluf3\ => \-aluf3\, aluf0a => aluf0a, aluf1a => aluf1a, aluf2a => aluf2a, aluf3a => aluf3a, yy1 => yy1, xx1 => xx1, yy0 => yy0, xx0 => xx0, \-cin32\ => \-cin32\, \-cin16\ => \-cin16\, \-cin0\ => \-cin0\, yout23 => yout23, xout23 => xout23, yout19 => yout19, xout19 => xout19, yout31 => yout31, xout31 => xout31, \-cin28\ => \-cin28\, \-cin24\ => \-cin24\, \-cin20\ => \-cin20\, yout27 => yout27, xout27 => xout27, yout7 => yout7, xout7 => xout7, yout3 => yout3, xout3 => xout3, yout15 => yout15, xout15 => xout15, \-cin12\ => \-cin12\, \-cin8\ => \-cin8\, \-cin4\ => \-cin4\, yout11 => yout11, xout11 => xout11, gnd => gnd, alusub => alusub, hi12 => hi12, \-ir3\ => \-ir3\, \-ir4\ => \-ir4\, aluadd => aluadd, ir6 => ir6, ir5 => ir5, ir7 => ir7, \-alumode\ => \-alumode\, \-ir2\ => \-ir2\, irjump => irjump, alumode => alumode, \-divposlasttime\ => \-divposlasttime\, q0 => q0, \-div\ => \-div\, divsubcond => divsubcond, divaddcond => divaddcond, a31b => a31b, \-a31\ => \-a31\, ir4 => ir4, ir3 => ir3, ir2 => ir2, \-ir1\ => \-ir1\, ir1 => ir1, \-ir0\ => \-ir0\, ir0 => ir0, a31a => a31a, \-mulnop\ => \-mulnop\, \-irjump\ => \-irjump\, \-mul\ => \-mul\, osel1a => osel1a, \-ir13\ => \-ir13\, \-iralu\ => \-iralu\, osel0a => osel0a, \-ir12\ => \-ir12\, osel1b => osel1b, osel0b => osel0b);
  i_alu0 : entity cadr_book.alu0(ttl) port map(a12 => a12, m12 => m12, aluf3b => aluf3b, aluf2b => aluf2b, aluf1b => aluf1b, aluf0b => aluf0b, \-cin12\ => \-cin12\, alumode => alumode, alu12 => alu12, alu13 => alu13, alu14 => alu14, alu15 => alu15, aeqm => aeqm, xout15 => xout15, yout15 => yout15, a15 => a15, m15 => m15, a14 => a14, m14 => m14, a13 => a13, m13 => m13, a4 => a4, m4 => m4, \-cin4\ => \-cin4\, alu4 => alu4, alu5 => alu5, alu6 => alu6, alu7 => alu7, xout7 => xout7, yout7 => yout7, a7 => a7, m7 => m7, a6 => a6, m6 => m6, a5 => a5, m5 => m5, a8 => a8, m8 => m8, \-cin8\ => \-cin8\, alu8 => alu8, alu9 => alu9, alu10 => alu10, alu11 => alu11, xout11 => xout11, yout11 => yout11, a11 => a11, m11 => m11, a10 => a10, m10 => m10, a9 => a9, m9 => m9, a0 => a0, m0 => m0, \-cin0\ => \-cin0\, alu0 => alu0, alu1 => alu1, alu2 => alu2, alu3 => alu3, xout3 => xout3, yout3 => yout3, a3 => a3, m3 => m3, a2 => a2, m2 => m2, a1 => a1, m1 => m1);
  i_alu1 : entity cadr_book.alu1(ttl) port map(a31a => a31a, m31b => m31b, aluf3a => aluf3a, aluf2a => aluf2a, aluf1a => aluf1a, aluf0a => aluf0a, \-cin32\ => \-cin32\, alumode => alumode, alu32 => alu32, m31 => m31, hi12 => hi12, a28 => a28, m28 => m28, \-cin28\ => \-cin28\, alu28 => alu28, alu29 => alu29, alu30 => alu30, alu31 => alu31, aeqm => aeqm, xout31 => xout31, yout31 => yout31, a31b => a31b, a30 => a30, m30 => m30, a29 => a29, m29 => m29, a20 => a20, m20 => m20, \-cin20\ => \-cin20\, alu20 => alu20, alu21 => alu21, alu22 => alu22, alu23 => alu23, xout23 => xout23, yout23 => yout23, a23 => a23, m23 => m23, a22 => a22, m22 => m22, a21 => a21, m21 => m21, a24 => a24, m24 => m24, \-cin24\ => \-cin24\, alu24 => alu24, alu25 => alu25, alu26 => alu26, alu27 => alu27, xout27 => xout27, yout27 => yout27, a27 => a27, m27 => m27, a26 => a26, m26 => m26, a25 => a25, m25 => m25, a16 => a16, m16 => m16, \-cin16\ => \-cin16\, alu16 => alu16, alu17 => alu17, alu18 => alu18, alu19 => alu19, xout19 => xout19, yout19 => yout19, a19 => a19, m19 => m19, a18 => a18, m18 => m18, a17 => a17, m17 => m17);


--- The Q Register (q)
  i_qctl : entity cadr_book.qctl(ttl) port map(\-qdrive\ => \-qdrive\, tse2 => tse2, srcq => srcq, q7 => q7, mf0 => mf0, q6 => q6, mf1 => mf1, q5 => q5, mf2 => mf2, q4 => q4, mf3 => mf3, q3 => q3, mf4 => mf4, q2 => q2, mf5 => mf5, q1 => q1, mf6 => mf6, q0 => q0, mf7 => mf7, qdrive => qdrive, q31 => q31, mf24 => mf24, q30 => q30, mf25 => mf25, q29 => q29, mf26 => mf26, q28 => q28, mf27 => mf27, q27 => q27, mf28 => mf28, q26 => q26, mf29 => mf29, q25 => q25, mf30 => mf30, q24 => q24, mf31 => mf31, q23 => q23, mf16 => mf16, q22 => q22, mf17 => mf17, q21 => q21, mf18 => mf18, q20 => q20, mf19 => mf19, q19 => q19, mf20 => mf20, q18 => q18, mf21 => mf21, q17 => q17, mf22 => mf22, q16 => q16, mf23 => mf23, q15 => q15, mf8 => mf8, q14 => q14, mf9 => mf9, q13 => q13, mf10 => mf10, q12 => q12, mf11 => mf11, q11 => q11, mf12 => mf12, q10 => q10, mf13 => mf13, q9 => q9, mf14 => mf14, q8 => q8, mf15 => mf15, \-srcq\ => \-srcq\, \-alu31\ => \-alu31\, alu31 => alu31, \-iralu\ => \-iralu\, \-ir1\ => \-ir1\, qs1 => qs1, \-ir0\ => \-ir0\, qs0 => qs0);
  i_q : entity cadr_book.q(ttl) port map(hi7 => hi7, q23 => q23, alu24 => alu24, alu25 => alu25, alu26 => alu26, alu27 => alu27, q28 => q28, qs0 => qs0, qs1 => qs1, clk2b => clk2b, q27 => q27, q26 => q26, q25 => q25, q24 => q24, alu28 => alu28, alu29 => alu29, alu30 => alu30, alu31 => alu31, alu0 => alu0, q31 => q31, q30 => q30, q29 => q29, q15 => q15, alu16 => alu16, alu17 => alu17, alu18 => alu18, alu19 => alu19, q20 => q20, q19 => q19, q18 => q18, q17 => q17, q16 => q16, alu20 => alu20, alu21 => alu21, alu22 => alu22, alu23 => alu23, q22 => q22, q21 => q21, q7 => q7, alu8 => alu8, alu9 => alu9, alu10 => alu10, alu11 => alu11, q12 => q12, q11 => q11, q10 => q10, q9 => q9, q8 => q8, alu12 => alu12, alu13 => alu13, alu14 => alu14, alu15 => alu15, q14 => q14, q13 => q13, \-alu31\ => \-alu31\, alu1 => alu1, alu2 => alu2, alu3 => alu3, q4 => q4, q3 => q3, q2 => q2, q1 => q1, q0 => q0, alu4 => alu4, alu5 => alu5, alu6 => alu6, alu7 => alu7, q6 => q6, q5 => q5);


--- The L Register (l)
  i_l : entity cadr_book.l(ttl) port map(gnd => gnd, l7 => l7, ob7 => ob7, ob6 => ob6, l6 => l6, l5 => l5, ob5 => ob5, ob4 => ob4, l4 => l4, clk3f => clk3f, l3 => l3, ob3 => ob3, ob2 => ob2, l2 => l2, l1 => l1, ob1 => ob1, ob0 => ob0, l0 => l0, l15 => l15, ob15 => ob15, ob14 => ob14, l14 => l14, l13 => l13, ob13 => ob13, ob12 => ob12, l12 => l12, l11 => l11, ob11 => ob11, ob10 => ob10, l10 => l10, l9 => l9, ob9 => ob9, ob8 => ob8, l8 => l8, l23 => l23, ob23 => ob23, ob22 => ob22, l22 => l22, l21 => l21, ob21 => ob21, ob20 => ob20, l20 => l20, l19 => l19, ob19 => ob19, ob18 => ob18, l18 => l18, l17 => l17, ob17 => ob17, ob16 => ob16, l16 => l16, l31 => l31, ob31 => ob31, ob30 => ob30, l30 => l30, l29 => l29, ob29 => ob29, ob28 => ob28, l28 => l28, l27 => l27, ob27 => ob27, ob26 => ob26, l26 => l26, l25 => l25, ob25 => ob25, ob24 => ob24, l24 => l24, lparl => lparl, \-lparm\ => \-lparm\, lparity => lparity, \-lparity\ => \-lparity\);


--- The Dispatch Memory (dsp)
  i_dspctl : entity cadr_book.dspctl(ttl) port map(dmask0 => dmask0, dmask1 => dmask1, dmask2 => dmask2, dmask3 => dmask3, dmask4 => dmask4, dmask5 => dmask5, dmask6 => dmask6, ir5 => ir5, ir6 => ir6, ir7 => ir7, gnd => gnd, \-irdisp\ => \-irdisp\, dc6 => dc6, ir38 => ir38, ir39 => ir39, dc7 => dc7, ir40 => ir40, dc8 => dc8, clk3e => clk3e, dc9 => dc9, ir41 => ir41, dc0 => dc0, ir32 => ir32, ir33 => ir33, dc1 => dc1, ir34 => ir34, dc2 => dc2, dc3 => dc3, ir35 => ir35, dc4 => dc4, ir36 => ir36, ir37 => ir37, dc5 => dc5, dpareven => dpareven, dispenb => dispenb, dparok => dparok, \-dparh\ => \-dparh\, dparl => dparl, hi4 => hi4, aa16 => aa16, aa17 => aa17, a17 => a17, a16 => a16, a15 => a15, aa8 => aa8, a14 => a14, aa9 => aa9, a13 => a13, aa10 => aa10, a12 => a12, aa11 => aa11, a11 => a11, aa12 => aa12, a10 => a10, aa13 => aa13, a9 => a9, aa14 => aa14, a8 => a8, aa15 => aa15, a7 => a7, aa0 => aa0, a6 => a6, aa1 => aa1, a5 => a5, aa2 => aa2, a4 => a4, aa3 => aa3, a3 => a3, aa4 => aa4, a2 => a2, aa5 => aa5, a1 => a1, aa6 => aa6, a0 => a0, aa7 => aa7, \-dmapbenb\ => \-dmapbenb\, ir8 => ir8, ir9 => ir9, dispwr => dispwr, \-funct2\ => \-funct2\, dpc9 => dpc9, dpc10 => dpc10, dpc11 => dpc11, dpc12 => dpc12, dpc13 => dpc13, dn => dn, dp => dp, dr => dr, dpar => dpar, dpc0 => dpc0, dpc1 => dpc1, dpc2 => dpc2, dpc3 => dpc3, dpc4 => dpc4, dpc5 => dpc5, dpc6 => dpc6, dpc7 => dpc7, dpc8 => dpc8);
  i_dram0 : entity cadr_book.dram0(ttl) port map(wp2 => wp2, dispwr => dispwr, \-dwea\ => \-dwea\, \-dadr10a\ => \-dadr10a\, dadr10a => dadr10a, ir22b => ir22b, \-dadr9a\ => \-dadr9a\, ir21b => ir21b, \-dadr8a\ => \-dadr8a\, ir20b => ir20b, \-dadr7a\ => \-dadr7a\, ir19b => ir19b, ir12b => ir12b, vmo19 => vmo19, ir9b => ir9b, r0 => r0, dmask0 => dmask0, \-dmapbenb\ => \-dmapbenb\, \-dadr0a\ => \-dadr0a\, vmo18 => vmo18, ir8b => ir8b, hi6 => hi6, gnd => gnd, ir12 => ir12, ir13 => ir13, ir18b => ir18b, ir14 => ir14, ir17b => ir17b, ir15 => ir15, ir16b => ir16b, ir16 => ir16, ir15b => ir15b, ir17 => ir17, ir14b => ir14b, ir18 => ir18, ir13b => ir13b, ir19 => ir19, \-dadr1a\ => \-dadr1a\, \-dadr2a\ => \-dadr2a\, \-dadr3a\ => \-dadr3a\, \-dadr4a\ => \-dadr4a\, dpc5 => dpc5, \-dadr5a\ => \-dadr5a\, \-dadr6a\ => \-dadr6a\, aa5 => aa5, dpc4 => dpc4, aa4 => aa4, r3 => r3, dmask6 => dmask6, r6 => r6, dmask3 => dmask3, dpc3 => dpc3, aa3 => aa3, dpc2 => dpc2, aa2 => aa2, r2 => r2, hi4 => hi4, dmask5 => dmask5, r5 => r5, dmask2 => dmask2, dpc1 => dpc1, aa1 => aa1, dpc0 => dpc0, aa0 => aa0, r1 => r1, dmask4 => dmask4, r4 => r4, dmask1 => dmask1);
  i_dram1 : entity cadr_book.dram1(ttl) port map(wp2 => wp2, dispwr => dispwr, \-dweb\ => \-dweb\, \-vmo19\ => \-vmo19\, vmo19 => vmo19, \-vmo18\ => \-vmo18\, vmo18 => vmo18, \-dadr9b\ => \-dadr9b\, ir21b => ir21b, \-dadr8b\ => \-dadr8b\, ir20b => ir20b, \-dadr7b\ => \-dadr7b\, ir19b => ir19b, ir12b => ir12b, ir9b => ir9b, r0 => r0, dmask0 => dmask0, \-dmapbenb\ => \-dmapbenb\, \-dadr0b\ => \-dadr0b\, ir8b => ir8b, hi6 => hi6, dadr10a => dadr10a, \-dadr1b\ => \-dadr1b\, \-dadr2b\ => \-dadr2b\, \-dadr3b\ => \-dadr3b\, \-dadr4b\ => \-dadr4b\, dpc11 => dpc11, \-dadr5b\ => \-dadr5b\, \-dadr6b\ => \-dadr6b\, aa11 => aa11, \-dadr10a\ => \-dadr10a\, dpc10 => dpc10, aa10 => aa10, r3 => r3, ir18b => ir18b, dmask6 => dmask6, r6 => r6, ir15b => ir15b, dmask3 => dmask3, dpc9 => dpc9, aa9 => aa9, dadr10c => dadr10c, dpc8 => dpc8, aa8 => aa8, \-dadr10c\ => \-dadr10c\, r2 => r2, ir17b => ir17b, dmask5 => dmask5, r5 => r5, ir14b => ir14b, dmask2 => dmask2, dpc7 => dpc7, aa7 => aa7, dpc6 => dpc6, aa6 => aa6, r1 => r1, ir16b => ir16b, dmask4 => dmask4, r4 => r4, ir13b => ir13b, dmask1 => dmask1, gnd => gnd, ir20 => ir20, ir21 => ir21, ir22 => ir22, ir8 => ir8, ir9 => ir9, ir22b => ir22b);
  i_dram2 : entity cadr_book.dram2(ttl) port map(dadr10c => dadr10c, \-dadr0c\ => \-dadr0c\, \-dadr1c\ => \-dadr1c\, \-dadr2c\ => \-dadr2c\, \-dadr3c\ => \-dadr3c\, \-dadr4c\ => \-dadr4c\, dpar => dpar, \-dadr5c\ => \-dadr5c\, \-dadr6c\ => \-dadr6c\, \-dadr7c\ => \-dadr7c\, \-dadr8c\ => \-dadr8c\, \-dadr9c\ => \-dadr9c\, \-dwec\ => \-dwec\, aa17 => aa17, \-dadr10c\ => \-dadr10c\, dr => dr, aa16 => aa16, r3 => r3, ir18b => ir18b, hi11 => hi11, dmask6 => dmask6, r6 => r6, ir15b => ir15b, dmask3 => dmask3, dp => dp, aa15 => aa15, dn => dn, aa14 => aa14, r2 => r2, ir17b => ir17b, dmask5 => dmask5, r5 => r5, ir14b => ir14b, dmask2 => dmask2, dpc13 => dpc13, aa13 => aa13, dpc12 => dpc12, aa12 => aa12, r1 => r1, ir16b => ir16b, dmask4 => dmask4, r4 => r4, ir13b => ir13b, dmask1 => dmask1, ir12b => ir12b, vmo19 => vmo19, ir9b => ir9b, r0 => r0, dmask0 => dmask0, \-dmapbenb\ => \-dmapbenb\, vmo18 => vmo18, ir8b => ir8b, hi6 => hi6, ir22b => ir22b, ir21b => ir21b, ir20b => ir20b, ir19b => ir19b, dispwr => dispwr, wp2 => wp2);


--- Jump Conditions (flag)
  i_flag : entity cadr_book.flag(ttl) port map(ir45 => ir45, \-nopa\ => \-nopa\, \-ilong\ => \-ilong\, ob29 => ob29, \lc_byte_mode\ => \lc_byte_mode\, ob28 => ob28, \prog.unibus.reset\ => \prog.unibus.reset\, hi4 => hi4, gnd => gnd, clk3c => clk3c, \int.enable\ => \int.enable\, ob27 => ob27, \sequence.break\ => \sequence.break\, ob26 => ob26, \-destintctl\ => \-destintctl\, \-reset\ => \-reset\, \-statbit\ => \-statbit\, ir46 => ir46, aeqm => aeqm, alu32 => alu32, aluneg => aluneg, r0 => r0, jcond => jcond, \-jcond\ => \-jcond\, conds2 => conds2, conds1 => conds1, conds0 => conds0, \pgf.or.int.or.sb\ => \pgf.or.int.or.sb\, \pgf.or.int\ => \pgf.or.int\, \-vmaok\ => \-vmaok\, ir2 => ir2, ir5 => ir5, ir1 => ir1, ir0 => ir0, \-alu32\ => \-alu32\, sint => sint, sintr => sintr);


--- Flow of Control (contrl)
  i_contrl : entity cadr_book.contrl(ttl) port map(spushd => spushd, tse3a => tse3a, spcwpass => spcwpass, \-ipopj\ => \-ipopj\, \-iwrited\ => \-iwrited\, \-popj\ => \-popj\, spcdrive => spcdrive, spcenb => spcenb, \-reset\ => \-reset\, inop => inop, \-inop\ => \-inop\, n => n, clk3c => clk3c, \-spushd\ => \-spushd\, spush => spush, iwrite => iwrite, iwrited => iwrited, \-srcspc\ => \-srcspc\, \-srcspcpop\ => \-srcspcpop\, \-spcdrive\ => \-spcdrive\, \-spcpass\ => \-spcpass\, \-spcwpass\ => \-spcwpass\, ir42 => ir42, \-nop\ => \-nop\, nop => nop, \-srcspcpopreal\ => \-srcspcpopreal\, \-nopa\ => \-nopa\, \-nop11\ => \-nop11\, \-irdisp\ => \-irdisp\, dr => dr, \-ignpopj\ => \-ignpopj\, \-destspc\ => \-destspc\, destspc => destspc, dp => dp, \-dfall\ => \-dfall\, \-trap\ => \-trap\, irdisp => irdisp, \-funct2\ => \-funct2\, dispenb => dispenb, irjump => irjump, ir6 => ir6, jfalse => jfalse, jcalf => jcalf, ir8 => ir8, jretf => jretf, jret => jret, ir7 => ir7, dn => dn, \-jcond\ => \-jcond\, hi4 => hi4, jcond => jcond, \-ir6\ => \-ir6\, \-dr\ => \-dr\, \-spush\ => \-spush\, pcs1 => pcs1, popj => popj, \-dp\ => \-dp\, \-spop\ => \-spop\, \-ir8\ => \-ir8\, ir9 => ir9, pcs0 => pcs0, \-spcnt\ => \-spcnt\, \-destspcd\ => \-destspcd\, destspcd => destspcd, wp4c => wp4c, \-swpb\ => \-swpb\, \-swpa\ => \-swpa\);


--- Microcode Subroutine Return Stack (spc)
  i_spc : entity cadr_book.spc(ttl) port map(\-swpa\ => \-swpa\, gnd => gnd, spcw14 => spcw14, spcptr4 => spcptr4, hi1 => hi1, spco14 => spco14, spco15 => spco15, spcptr3 => spcptr3, spcptr2 => spcptr2, spcptr1 => spcptr1, spcptr0 => spcptr0, spcw15 => spcw15, spcw12 => spcw12, spco12 => spco12, spco13 => spco13, spcw13 => spcw13, spcw10 => spcw10, spco10 => spco10, spco11 => spco11, spcw11 => spcw11, spcopar => spcopar, spco18 => spco18, spco17 => spco17, spco16 => spco16, hi2 => hi2, hi3 => hi3, hi4 => hi4, hi5 => hi5, hi6 => hi6, hi7 => hi7, \-swpb\ => \-swpb\, spcw4 => spcw4, spco4 => spco4, spco5 => spco5, spcw5 => spcw5, spcw2 => spcw2, spco2 => spco2, spco3 => spco3, spcw3 => spcw3, spcw0 => spcw0, spco0 => spco0, spco1 => spco1, spcw1 => spcw1, spco9 => spco9, spco8 => spco8, spco7 => spco7, spco6 => spco6, hi8 => hi8, hi9 => hi9, hi10 => hi10, hi11 => hi11, hi12 => hi12, spush => spush, clk4f => clk4f, \-spcnt\ => \-spcnt\, \-spccry\ => \-spccry\, spcw18 => spcw18, spcwpar => spcwpar, spcw16 => spcw16, spcw17 => spcw17, spcw8 => spcw8, spcw9 => spcw9, spcw6 => spcw6, spcw7 => spcw7);
  i_spclch : entity cadr_book.spclch(ttl) port map(\-spcdrive\ => \-spcdrive\, m23 => m23, gnd => gnd, m22 => m22, m21 => m21, m20 => m20, clk4c => clk4c, m19 => m19, spco18 => spco18, m18 => m18, m17 => m17, spco17 => spco17, spco16 => spco16, m16 => m16, m15 => m15, spco15 => spco15, spco14 => spco14, m14 => m14, m13 => m13, spco13 => spco13, spco12 => spco12, m12 => m12, m11 => m11, spco11 => spco11, spco10 => spco10, m10 => m10, m9 => m9, spco9 => spco9, spco8 => spco8, m8 => m8, m7 => m7, spco7 => spco7, spco6 => spco6, m6 => m6, m5 => m5, spco5 => spco5, spco4 => spco4, m4 => m4, m3 => m3, spco3 => spco3, spco2 => spco2, m2 => m2, m1 => m1, spco1 => spco1, spco0 => spco0, m0 => m0, m24 => m24, m25 => m25, m26 => m26, spcptr4 => spcptr4, m27 => m27, spcptr3 => spcptr3, m28 => m28, spcptr2 => spcptr2, m29 => m29, spcptr1 => spcptr1, m30 => m30, spcptr0 => spcptr0, m31 => m31, spcdrive => spcdrive, hi1 => hi1, spc16 => spc16, spc17 => spc17, spc18 => spc18, spcpar => spcpar, spcwpar => spcwpar, spcw18 => spcw18, spcw17 => spcw17, spcw16 => spcw16, spcwpass => spcwpass, \-spcwpass\ => \-spcwpass\, spcw15 => spcw15, spc8 => spc8, spcw14 => spcw14, spc9 => spc9, spcw13 => spcw13, spc10 => spc10, spcw12 => spcw12, spc11 => spc11, spcw11 => spcw11, spc12 => spc12, spcw10 => spcw10, spc13 => spc13, spcw9 => spcw9, spc14 => spc14, spcw8 => spcw8, spc15 => spc15, spcw7 => spcw7, spc0 => spc0, spcw6 => spcw6, spc1 => spc1, spcw5 => spcw5, spc2 => spc2, spcw4 => spcw4, spc3 => spc3, spcw3 => spcw3, spc4 => spc4, spcw2 => spcw2, spc5 => spc5, spcw1 => spcw1, spc6 => spc6, spcw0 => spcw0, spc7 => spc7, \-spcpass\ => \-spcpass\, clk4d => clk4d, spcopar => spcopar);
  i_spcw : entity cadr_book.spcw(ttl) port map(destspcd => destspcd, reta12 => reta12, l12 => l12, spcw12 => spcw12, reta13 => reta13, l13 => l13, spcw13 => spcw13, spcw14 => spcw14, l14 => l14, gnd => gnd, spcw15 => spcw15, l15 => l15, reta8 => reta8, l8 => l8, spcw8 => spcw8, reta9 => reta9, l9 => l9, spcw9 => spcw9, spcw10 => spcw10, l10 => l10, reta10 => reta10, spcw11 => spcw11, l11 => l11, reta11 => reta11, reta4 => reta4, l4 => l4, spcw4 => spcw4, reta5 => reta5, l5 => l5, spcw5 => spcw5, spcw6 => spcw6, l6 => l6, reta6 => reta6, spcw7 => spcw7, l7 => l7, reta7 => reta7, reta0 => reta0, l0 => l0, spcw0 => spcw0, reta1 => reta1, l1 => l1, spcw1 => spcw1, spcw2 => spcw2, l2 => l2, reta2 => reta2, spcw3 => spcw3, l3 => l3, reta3 => reta3, n => n, ipc12 => ipc12, wpc12 => wpc12, wpc13 => wpc13, ipc13 => ipc13, clk4d => clk4d, ipc8 => ipc8, wpc8 => wpc8, wpc9 => wpc9, ipc9 => ipc9, ipc10 => ipc10, wpc10 => wpc10, wpc11 => wpc11, ipc11 => ipc11, ipc4 => ipc4, wpc4 => wpc4, wpc5 => wpc5, ipc5 => ipc5, ipc6 => ipc6, wpc6 => wpc6, wpc7 => wpc7, ipc7 => ipc7, ipc0 => ipc0, wpc0 => wpc0, wpc1 => wpc1, ipc1 => ipc1, ipc2 => ipc2, wpc2 => wpc2, wpc3 => wpc3, ipc3 => ipc3, l16 => l16, spcw16 => spcw16, l17 => l17, spcw17 => spcw17, spcw18 => spcw18, l18 => l18);
  i_spcpar : entity cadr_book.spcpar(ttl) port map(spcwparh => spcwparh, \-spcwparl\ => \-spcwparl\, spcwpar => spcwpar, spcw17 => spcw17, spcw18 => spcw18, gnd => gnd, spcw12 => spcw12, spcw13 => spcw13, spcw14 => spcw14, spcw15 => spcw15, spcw16 => spcw16, spcw5 => spcw5, spcw6 => spcw6, spcw7 => spcw7, spcw8 => spcw8, spcw9 => spcw9, spcw10 => spcw10, spcw11 => spcw11, spcw0 => spcw0, spcw1 => spcw1, spcw2 => spcw2, spcw3 => spcw3, spcw4 => spcw4, spc16 => spc16, spc17 => spc17, spc18 => spc18, spcpar => spcpar, spcparh => spcparh, spc11 => spc11, spc12 => spc12, spc13 => spc13, spc14 => spc14, spc15 => spc15, spc5 => spc5, spc6 => spc6, spc7 => spc7, spc8 => spc8, spc9 => spc9, spc10 => spc10, spcparok => spcparok, spc0 => spc0, spc1 => spc1, spc2 => spc2, spc3 => spc3, spc4 => spc4);
  i_lpc : entity cadr_book.lpc(ttl) port map(gnd => gnd, pc8 => pc8, pc9 => pc9, pc10 => pc10, pc13b => pc13b, pc11 => pc11, pc12b => pc12b, pc12 => pc12, pc11b => pc11b, pc13 => pc13, pc10b => pc10b, pc9b => pc9b, pc8b => pc8b, hi5 => hi5, pc0 => pc0, pc7b => pc7b, pc1 => pc1, pc6b => pc6b, pc2 => pc2, pc5b => pc5b, pc3 => pc3, pc4b => pc4b, pc4 => pc4, pc3b => pc3b, pc5 => pc5, pc2b => pc2b, pc6 => pc6, pc1b => pc1b, pc7 => pc7, pc0b => pc0b, irdisp => irdisp, ir25 => ir25, lpc12 => lpc12, wpc12 => wpc12, lpc13 => lpc13, wpc13 => wpc13, lpc8 => lpc8, wpc8 => wpc8, lpc9 => lpc9, wpc9 => wpc9, wpc10 => wpc10, lpc10 => lpc10, wpc11 => wpc11, lpc11 => lpc11, lpc4 => lpc4, wpc4 => wpc4, lpc5 => lpc5, wpc5 => wpc5, wpc6 => wpc6, lpc6 => lpc6, wpc7 => wpc7, lpc7 => lpc7, lpc0 => lpc0, wpc0 => wpc0, lpc1 => lpc1, wpc1 => wpc1, wpc2 => wpc2, lpc2 => lpc2, wpc3 => wpc3, lpc3 => lpc3, \lpc.hold\ => \lpc.hold\, clk4b => clk4b);


--- Next PC Selector (npc)
  i_npc : entity cadr_book.npc(ttl) port map(ipc13 => ipc13, gnd => gnd, pc13 => pc13, ipc12 => ipc12, pc12 => pc12, pccry11 => pccry11, ipc9 => ipc9, pc9 => pc9, ipc8 => ipc8, pc8 => pc8, pccry7 => pccry7, ipc11 => ipc11, pc11 => pc11, ipc10 => ipc10, pc10 => pc10, ipc5 => ipc5, pc5 => pc5, ipc4 => ipc4, pc4 => pc4, pccry3 => pccry3, ipc7 => ipc7, pc7 => pc7, ipc6 => ipc6, pc6 => pc6, ipc1 => ipc1, pc1 => pc1, ipc0 => ipc0, pc0 => pc0, hi4 => hi4, ipc3 => ipc3, pc3 => pc3, ipc2 => ipc2, pc2 => pc2, trapb => trapb, pcs1 => pcs1, dpc3 => dpc3, ir15 => ir15, spc3 => spc3, npc3 => npc3, npc2 => npc2, spc2 => spc2, ir14 => ir14, dpc2 => dpc2, pcs0 => pcs0, dpc1 => dpc1, ir13 => ir13, spc1a => spc1a, npc1 => npc1, npc0 => npc0, spc0 => spc0, ir12 => ir12, dpc0 => dpc0, npc13 => npc13, npc12 => npc12, clk4b => clk4b, npc11 => npc11, npc10 => npc10, npc9 => npc9, npc8 => npc8, npc7 => npc7, npc6 => npc6, npc5 => npc5, npc4 => npc4, trapa => trapa, dpc13 => dpc13, ir25 => ir25, spc13 => spc13, spc12 => spc12, ir24 => ir24, dpc12 => dpc12, dpc11 => dpc11, ir23 => ir23, spc11 => spc11, spc10 => spc10, ir22 => ir22, dpc10 => dpc10, dpc9 => dpc9, ir21 => ir21, spc9 => spc9, spc8 => spc8, ir20 => ir20, dpc8 => dpc8, dpc7 => dpc7, ir19 => ir19, spc7 => spc7, spc6 => spc6, ir18 => ir18, dpc6 => dpc6, dpc5 => dpc5, ir17 => ir17, spc5 => spc5, spc4 => spc4, ir16 => ir16, dpc4 => dpc4);


--- The LC register and Instruction Prefetch (lc)
  i_lc : entity cadr_book.lc(ttl) port map(\-lcdrive\ => \-lcdrive\, needfetch => needfetch, mf24 => mf24, gnd => gnd, mf25 => mf25, \lc_byte_mode\ => \lc_byte_mode\, mf26 => mf26, \prog.unibus.reset\ => \prog.unibus.reset\, mf27 => mf27, \int.enable\ => \int.enable\, mf28 => mf28, \sequence.break\ => \sequence.break\, mf29 => mf29, lc25 => lc25, mf30 => mf30, lc24 => lc24, mf31 => mf31, lcdrive => lcdrive, srclc => srclc, tse1a => tse1a, lc7 => lc7, mf0 => mf0, lc6 => lc6, mf1 => mf1, lc5 => lc5, mf2 => mf2, lc4 => lc4, mf3 => mf3, lc3 => lc3, mf4 => mf4, lc2 => lc2, mf5 => mf5, lc1 => lc1, mf6 => mf6, lc0b => lc0b, mf7 => mf7, lc23 => lc23, mf16 => mf16, lc22 => lc22, mf17 => mf17, lc21 => lc21, mf18 => mf18, lc20 => lc20, mf19 => mf19, lc19 => lc19, mf20 => mf20, lc18 => lc18, mf21 => mf21, lc17 => lc17, mf22 => mf22, lc16 => lc16, mf23 => mf23, lc15 => lc15, mf8 => mf8, lc14 => lc14, mf9 => mf9, lc13 => lc13, mf10 => mf10, lc12 => lc12, mf11 => mf11, lc11 => lc11, mf12 => mf12, lc10 => lc10, mf13 => mf13, lc9 => lc9, mf14 => mf14, lc8 => lc8, mf15 => mf15, hi11 => hi11, clk1a => clk1a, ob20 => ob20, ob21 => ob21, ob22 => ob22, ob23 => ob23, \-destlc\ => \-destlc\, \-lcry19\ => \-lcry19\, \-lcry23\ => \-lcry23\, ob16 => ob16, ob17 => ob17, ob18 => ob18, ob19 => ob19, \-lcry15\ => \-lcry15\, clk2a => clk2a, ob12 => ob12, ob13 => ob13, ob14 => ob14, ob15 => ob15, \-lcry11\ => \-lcry11\, clk2c => clk2c, ob8 => ob8, ob9 => ob9, ob10 => ob10, ob11 => ob11, \-lcry7\ => \-lcry7\, \-srclc\ => \-srclc\, ob24 => ob24, ob25 => ob25, ob4 => ob4, ob5 => ob5, ob6 => ob6, ob7 => ob7, \-lcry3\ => \-lcry3\);
  i_lcc : entity cadr_book.lcc(ttl) port map(\lc_byte_mode\ => \lc_byte_mode\, \-lcinc\ => \-lcinc\, lca1 => lca1, gnd => gnd, lc1 => lc1, lca0 => lca0, lc0 => lc0, lcinc => lcinc, lcry3 => lcry3, lca3 => lca3, lc3 => lc3, lca2 => lca2, lc2 => lc2, \-destlc\ => \-destlc\, ob3 => ob3, ob2 => ob2, clk2a => clk2a, ob1 => ob1, ob0 => ob0, lc0b => lc0b, \inst_in_left_half\ => \inst_in_left_half\, \-ir4\ => \-ir4\, \-sh4\ => \-sh4\, \-sh3\ => \-sh3\, \-ir3\ => \-ir3\, \inst_in_2nd_or_4th_quarter\ => \inst_in_2nd_or_4th_quarter\, \-lc_modifies_mrot\ => \-lc_modifies_mrot\, spc14 => spc14, \-srcspcpopreal\ => \-srcspcpopreal\, \-ifetch\ => \-ifetch\, needfetch => needfetch, \have_wrong_word\ => \have_wrong_word\, \last_byte_in_word\ => \last_byte_in_word\, ir10 => ir10, ir11 => ir11, \-newlc\ => \-newlc\, \-newlc.in\ => \-newlc.in\, \-reset\ => \-reset\, newlc => newlc, int => int, sintr => sintr, clk3c => clk3c, \next.instrd\ => \next.instrd\, \next.instr\ => \next.instr\, \-spop\ => \-spop\, \-needfetch\ => \-needfetch\, spcmung => spcmung, ir24 => ir24, irdisp => irdisp, spc1 => spc1, spc1a => spc1a);


--- The VMA and VMA Selector (vma)
  i_vma : entity cadr_book.vma(ttl) port map(\-vmadrive\ => \-vmadrive\, \-vma31\ => \-vma31\, mf24 => mf24, \-vma30\ => \-vma30\, mf25 => mf25, \-vma29\ => \-vma29\, mf26 => mf26, \-vma28\ => \-vma28\, mf27 => mf27, \-vma27\ => \-vma27\, mf28 => mf28, \-vma26\ => \-vma26\, mf29 => mf29, \-vma25\ => \-vma25\, mf30 => mf30, \-vma24\ => \-vma24\, mf31 => mf31, \-vma7\ => \-vma7\, mf0 => mf0, \-vma6\ => \-vma6\, mf1 => mf1, \-vma5\ => \-vma5\, mf2 => mf2, \-vma4\ => \-vma4\, mf3 => mf3, \-vma3\ => \-vma3\, mf4 => mf4, \-vma2\ => \-vma2\, mf5 => mf5, \-vma1\ => \-vma1\, mf6 => mf6, \-vma0\ => \-vma0\, mf7 => mf7, \-vma23\ => \-vma23\, mf16 => mf16, \-vma22\ => \-vma22\, mf17 => mf17, \-vma21\ => \-vma21\, mf18 => mf18, \-vma20\ => \-vma20\, mf19 => mf19, \-vma19\ => \-vma19\, mf20 => mf20, \-vma18\ => \-vma18\, mf21 => mf21, \-vma17\ => \-vma17\, mf22 => mf22, \-vma16\ => \-vma16\, mf23 => mf23, \-vma15\ => \-vma15\, mf8 => mf8, \-vma14\ => \-vma14\, mf9 => mf9, \-vma13\ => \-vma13\, mf10 => mf10, \-vma12\ => \-vma12\, mf11 => mf11, \-vma11\ => \-vma11\, mf12 => mf12, \-vma10\ => \-vma10\, mf13 => mf13, \-vma9\ => \-vma9\, mf14 => mf14, \-vma8\ => \-vma8\, mf15 => mf15, tse2 => tse2, srcvma => srcvma, \-vmaenb\ => \-vmaenb\, \-vmas24\ => \-vmas24\, \-vmas25\ => \-vmas25\, \-vmas26\ => \-vmas26\, clk1a => clk1a, \-vmas27\ => \-vmas27\, \-vmas28\ => \-vmas28\, \-vmas29\ => \-vmas29\, \-vmas30\ => \-vmas30\, \-vmas31\ => \-vmas31\, \-vmas0\ => \-vmas0\, \-vmas1\ => \-vmas1\, \-vmas2\ => \-vmas2\, clk2a => clk2a, \-vmas3\ => \-vmas3\, \-vmas4\ => \-vmas4\, \-vmas5\ => \-vmas5\, \-vmas12\ => \-vmas12\, \-vmas13\ => \-vmas13\, \-vmas14\ => \-vmas14\, \-vmas15\ => \-vmas15\, \-vmas16\ => \-vmas16\, \-vmas17\ => \-vmas17\, \-vmas18\ => \-vmas18\, \-vmas19\ => \-vmas19\, \-vmas20\ => \-vmas20\, \-vmas21\ => \-vmas21\, \-vmas22\ => \-vmas22\, \-vmas23\ => \-vmas23\, \-vmas6\ => \-vmas6\, \-vmas7\ => \-vmas7\, \-vmas8\ => \-vmas8\, clk2c => clk2c, \-vmas9\ => \-vmas9\, \-vmas10\ => \-vmas10\, \-vmas11\ => \-vmas11\, \-srcvma\ => \-srcvma\);
  i_vmas : entity cadr_book.vmas(ttl) port map(vmasela => vmasela, lc22 => lc22, ob20 => ob20, \-vmas20\ => \-vmas20\, lc23 => lc23, ob21 => ob21, \-vmas21\ => \-vmas21\, \-vmas22\ => \-vmas22\, ob22 => ob22, lc24 => lc24, \-vmas23\ => \-vmas23\, ob23 => ob23, lc25 => lc25, gnd => gnd, ob28 => ob28, \-vmas28\ => \-vmas28\, ob29 => ob29, \-vmas29\ => \-vmas29\, \-vmas30\ => \-vmas30\, ob30 => ob30, \-vmas31\ => \-vmas31\, ob31 => ob31, vmaselb => vmaselb, lc14 => lc14, ob12 => ob12, \-vmas12\ => \-vmas12\, lc15 => lc15, ob13 => ob13, \-vmas13\ => \-vmas13\, \-vmas14\ => \-vmas14\, ob14 => ob14, lc16 => lc16, \-vmas15\ => \-vmas15\, ob15 => ob15, lc17 => lc17, lc18 => lc18, ob16 => ob16, \-vmas16\ => \-vmas16\, lc19 => lc19, ob17 => ob17, \-vmas17\ => \-vmas17\, \-vmas18\ => \-vmas18\, ob18 => ob18, lc20 => lc20, \-vmas19\ => \-vmas19\, ob19 => ob19, lc21 => lc21, \-memstart\ => \-memstart\, \-vma12\ => \-vma12\, \-md12\ => \-md12\, mapi12 => mapi12, \-vma13\ => \-vma13\, \-md13\ => \-md13\, mapi13 => mapi13, mapi14 => mapi14, \-md14\ => \-md14\, \-vma14\ => \-vma14\, mapi15 => mapi15, \-md15\ => \-md15\, \-vma15\ => \-vma15\, \-vma16\ => \-vma16\, \-md16\ => \-md16\, mapi16 => mapi16, \-vma17\ => \-vma17\, \-md17\ => \-md17\, mapi17 => mapi17, mapi18 => mapi18, \-md18\ => \-md18\, \-vma18\ => \-vma18\, mapi19 => mapi19, \-md19\ => \-md19\, \-vma19\ => \-vma19\, \-vma20\ => \-vma20\, \-md20\ => \-md20\, mapi20 => mapi20, \-vma21\ => \-vma21\, \-md21\ => \-md21\, mapi21 => mapi21, mapi22 => mapi22, \-md22\ => \-md22\, \-vma22\ => \-vma22\, mapi23 => mapi23, \-md23\ => \-md23\, \-vma23\ => \-vma23\, lc2 => lc2, ob0 => ob0, \-vmas0\ => \-vmas0\, lc3 => lc3, ob1 => ob1, \-vmas1\ => \-vmas1\, \-vmas2\ => \-vmas2\, ob2 => ob2, lc4 => lc4, \-vmas3\ => \-vmas3\, ob3 => ob3, lc5 => lc5, \-vma8\ => \-vma8\, \-md8\ => \-md8\, mapi8 => mapi8, \-vma9\ => \-vma9\, \-md9\ => \-md9\, mapi9 => mapi9, mapi10 => mapi10, \-md10\ => \-md10\, \-vma10\ => \-vma10\, mapi11 => mapi11, \-md11\ => \-md11\, \-vma11\ => \-vma11\, lc10 => lc10, ob8 => ob8, \-vmas8\ => \-vmas8\, lc11 => lc11, ob9 => ob9, \-vmas9\ => \-vmas9\, \-vmas10\ => \-vmas10\, ob10 => ob10, lc12 => lc12, \-vmas11\ => \-vmas11\, ob11 => ob11, lc13 => lc13, lc6 => lc6, ob4 => ob4, \-vmas4\ => \-vmas4\, lc7 => lc7, ob5 => ob5, \-vmas5\ => \-vmas5\, \-vmas6\ => \-vmas6\, ob6 => ob6, lc8 => lc8, \-vmas7\ => \-vmas7\, ob7 => ob7, lc9 => lc9, ob24 => ob24, \-vmas24\ => \-vmas24\, ob25 => ob25, \-vmas25\ => \-vmas25\, \-vmas26\ => \-vmas26\, ob26 => ob26, \-vmas27\ => \-vmas27\, ob27 => ob27);


--- The MD and the MD Selector (md)
  i_md : entity cadr_book.md(ttl) port map(\-mddrive\ => \-mddrive\, \-md31\ => \-md31\, mf24 => mf24, \-md30\ => \-md30\, mf25 => mf25, \-md29\ => \-md29\, mf26 => mf26, \-md28\ => \-md28\, mf27 => mf27, \-md27\ => \-md27\, mf28 => mf28, \-md26\ => \-md26\, mf29 => mf29, \-md25\ => \-md25\, mf30 => mf30, \-md24\ => \-md24\, mf31 => mf31, \-md23\ => \-md23\, mf16 => mf16, \-md22\ => \-md22\, mf17 => mf17, \-md21\ => \-md21\, mf18 => mf18, \-md20\ => \-md20\, mf19 => mf19, \-md19\ => \-md19\, mf20 => mf20, \-md18\ => \-md18\, mf21 => mf21, \-md17\ => \-md17\, mf22 => mf22, \-md16\ => \-md16\, mf23 => mf23, \-md7\ => \-md7\, mf0 => mf0, \-md6\ => \-md6\, mf1 => mf1, \-md5\ => \-md5\, mf2 => mf2, \-md4\ => \-md4\, mf3 => mf3, \-md3\ => \-md3\, mf4 => mf4, \-md2\ => \-md2\, mf5 => mf5, \-md1\ => \-md1\, mf6 => mf6, \-md0\ => \-md0\, mf7 => mf7, srcmd => srcmd, tse2 => tse2, \-md15\ => \-md15\, mf8 => mf8, \-md14\ => \-md14\, mf9 => mf9, \-md13\ => \-md13\, mf10 => mf10, \-md12\ => \-md12\, mf11 => mf11, \-md11\ => \-md11\, mf12 => mf12, \-md10\ => \-md10\, mf13 => mf13, \-md9\ => \-md9\, mf14 => mf14, \-md8\ => \-md8\, mf15 => mf15, gnd => gnd, \-mds31\ => \-mds31\, \-mds30\ => \-mds30\, \-mds29\ => \-mds29\, \-mds28\ => \-mds28\, mdclk => mdclk, \-mds27\ => \-mds27\, \-mds26\ => \-mds26\, \-mds25\ => \-mds25\, \-mds24\ => \-mds24\, \-mds7\ => \-mds7\, \-mds6\ => \-mds6\, \-mds5\ => \-mds5\, \-mds4\ => \-mds4\, \-mds3\ => \-mds3\, \-mds2\ => \-mds2\, \-mds1\ => \-mds1\, \-mds0\ => \-mds0\, \-mds23\ => \-mds23\, \-mds22\ => \-mds22\, \-mds21\ => \-mds21\, \-mds20\ => \-mds20\, \-mds19\ => \-mds19\, \-mds18\ => \-mds18\, \-mds17\ => \-mds17\, \-mds16\ => \-mds16\, destmdr => destmdr, \-clk2c\ => \-clk2c\, loadmd => loadmd, \-loadmd\ => \-loadmd\, \-destmdr\ => \-destmdr\, \-mds15\ => \-mds15\, \-mds14\ => \-mds14\, \-mds13\ => \-mds13\, \-mds12\ => \-mds12\, \-mds11\ => \-mds11\, \-mds10\ => \-mds10\, \-mds9\ => \-mds9\, \-mds8\ => \-mds8\, mdgetspar => mdgetspar, \-ignpar\ => \-ignpar\, mdhaspar => mdhaspar, \mempar_in\ => \mempar_in\, mdpar => mdpar, \-srcmd\ => \-srcmd\);
  i_mds : entity cadr_book.mds(ttl) port map(\-memdrive.a\ => \-memdrive.a\, \-md31\ => \-md31\, mem24 => mem24, \-md30\ => \-md30\, mem25 => mem25, \-md29\ => \-md29\, mem26 => mem26, \-md28\ => \-md28\, mem27 => mem27, \-md27\ => \-md27\, mem28 => mem28, \-md26\ => \-md26\, mem29 => mem29, \-md25\ => \-md25\, mem30 => mem30, \-md24\ => \-md24\, mem31 => mem31, \-memdrive.b\ => \-memdrive.b\, \-md7\ => \-md7\, mem0 => mem0, \-md6\ => \-md6\, mem1 => mem1, \-md5\ => \-md5\, mem2 => mem2, \-md4\ => \-md4\, mem3 => mem3, \-md3\ => \-md3\, mem4 => mem4, \-md2\ => \-md2\, mem5 => mem5, \-md1\ => \-md1\, mem6 => mem6, \-md0\ => \-md0\, mem7 => mem7, \-md23\ => \-md23\, mem16 => mem16, \-md22\ => \-md22\, mem17 => mem17, \-md21\ => \-md21\, mem18 => mem18, \-md20\ => \-md20\, mem19 => mem19, \-md19\ => \-md19\, mem20 => mem20, \-md18\ => \-md18\, mem21 => mem21, \-md17\ => \-md17\, mem22 => mem22, \-md16\ => \-md16\, mem23 => mem23, \-md15\ => \-md15\, mem8 => mem8, \-md14\ => \-md14\, mem9 => mem9, \-md13\ => \-md13\, mem10 => mem10, \-md12\ => \-md12\, mem11 => mem11, \-md11\ => \-md11\, mem12 => mem12, \-md10\ => \-md10\, mem13 => mem13, \-md9\ => \-md9\, mem14 => mem14, \-md8\ => \-md8\, mem15 => mem15, mdsela => mdsela, ob20 => ob20, \-mds20\ => \-mds20\, ob21 => ob21, \-mds21\ => \-mds21\, \-mds22\ => \-mds22\, ob22 => ob22, \-mds23\ => \-mds23\, ob23 => ob23, gnd => gnd, ob28 => ob28, \-mds28\ => \-mds28\, ob29 => ob29, \-mds29\ => \-mds29\, \-mds30\ => \-mds30\, ob30 => ob30, \-mds31\ => \-mds31\, ob31 => ob31, mdparodd => mdparodd, \mempar_out\ => \mempar_out\, hi11 => hi11, mdselb => mdselb, ob12 => ob12, \-mds12\ => \-mds12\, ob13 => ob13, \-mds13\ => \-mds13\, \-mds14\ => \-mds14\, ob14 => ob14, \-mds15\ => \-mds15\, ob15 => ob15, ob16 => ob16, \-mds16\ => \-mds16\, ob17 => ob17, \-mds17\ => \-mds17\, \-mds18\ => \-mds18\, ob18 => ob18, \-mds19\ => \-mds19\, ob19 => ob19, ob8 => ob8, \-mds8\ => \-mds8\, ob9 => ob9, \-mds9\ => \-mds9\, \-mds10\ => \-mds10\, ob10 => ob10, \-mds11\ => \-mds11\, ob11 => ob11, ob0 => ob0, \-mds0\ => \-mds0\, ob1 => ob1, \-mds1\ => \-mds1\, \-mds2\ => \-mds2\, ob2 => ob2, \-mds3\ => \-mds3\, ob3 => ob3, ob4 => ob4, \-mds4\ => \-mds4\, ob5 => ob5, \-mds5\ => \-mds5\, \-mds6\ => \-mds6\, ob6 => ob6, \-mds7\ => \-mds7\, ob7 => ob7, ob24 => ob24, \-mds24\ => \-mds24\, ob25 => ob25, \-mds25\ => \-mds25\, \-mds26\ => \-mds26\, ob26 => ob26, \-mds27\ => \-mds27\, ob27 => ob27);


--- First and Second Level Maps (vmem)
  i_vmem0 : entity cadr_book.vmem0(ttl) port map(\-vmap0\ => \-vmap0\, \-vmap1\ => \-vmap1\, \-vmap2\ => \-vmap2\, \-vmap3\ => \-vmap3\, \-vmap4\ => \-vmap4\, vpari => vpari, gnd => gnd, \-vma27\ => \-vma27\, \-vma28\ => \-vma28\, \-vma29\ => \-vma29\, vm0pari => vm0pari, \-vma30\ => \-vma30\, \-vma31\ => \-vma31\, \-mapi23\ => \-mapi23\, mapi22 => mapi22, mapi21 => mapi21, mapi20 => mapi20, mapi19 => mapi19, mapi18 => mapi18, mapi17 => mapi17, mapi16 => mapi16, mapi15 => mapi15, mapi14 => mapi14, mapi13 => mapi13, \-vm0wpb\ => \-vm0wpb\, mapi23 => mapi23, \-vm0wpa\ => \-vm0wpa\, memstart => memstart, srcmap => srcmap, \-use.map\ => \-use.map\, v0parok => v0parok, vmoparodd => vmoparodd, vmoparok => vmoparok);
  i_vmem1 : entity cadr_book.vmem1(ttl) port map(\-vma17\ => \-vma17\, \-vma18\ => \-vma18\, \-vma19\ => \-vma19\, \-vma20\ => \-vma20\, \-vma21\ => \-vma21\, \-vma22\ => \-vma22\, \-vma23\ => \-vma23\, vm1mpar => vm1mpar, \-vma12\ => \-vma12\, \-vma13\ => \-vma13\, \-vma14\ => \-vma14\, \-vma15\ => \-vma15\, \-vma16\ => \-vma16\, \-vma5\ => \-vma5\, \-vma6\ => \-vma6\, \-vma7\ => \-vma7\, \-vma8\ => \-vma8\, \-vma9\ => \-vma9\, \-vma10\ => \-vma10\, \-vma11\ => \-vma11\, \-vm1lpar\ => \-vm1lpar\, \-vma0\ => \-vma0\, \-vma1\ => \-vma1\, \-vma2\ => \-vma2\, \-vma3\ => \-vma3\, \-vma4\ => \-vma4\, gnd => gnd, vmap4a => vmap4a, vmap3a => vmap3a, vmap2a => vmap2a, vmap1a => vmap1a, vmap0a => vmap0a, \-vmo10\ => \-vmo10\, \-mapi12a\ => \-mapi12a\, \-mapi11a\ => \-mapi11a\, \-mapi10a\ => \-mapi10a\, \-mapi9a\ => \-mapi9a\, \-mapi8a\ => \-mapi8a\, \-vm1wpa\ => \-vm1wpa\, \-vmo4\ => \-vmo4\, \-vmo2\ => \-vmo2\, mapi10 => mapi10, mapi9 => mapi9, mapi8 => mapi8, \-vmap4\ => \-vmap4\, \-vmap3\ => \-vmap3\, \-vmap2\ => \-vmap2\, \-vmap1\ => \-vmap1\, \-vmap0\ => \-vmap0\, \-vmo0\ => \-vmo0\, vm1pari => vm1pari, mapi12 => mapi12, mapi11 => mapi11, \-mapi8b\ => \-mapi8b\, \-mapi9b\ => \-mapi9b\, \-mapi10b\ => \-mapi10b\, \-mapi11b\ => \-mapi11b\, \-mapi12b\ => \-mapi12b\, \-vmo11\ => \-vmo11\, \-vmo5\ => \-vmo5\, \-vmo9\ => \-vmo9\, \-vmo3\ => \-vmo3\, \-vmo8\ => \-vmo8\, \-vmo7\ => \-vmo7\, \-vmo1\ => \-vmo1\, \-vmo6\ => \-vmo6\);
  i_vmem2 : entity cadr_book.vmem2(ttl) port map(gnd => gnd, vmap4b => vmap4b, vmap3b => vmap3b, vmap2b => vmap2b, vmap1b => vmap1b, vmap0b => vmap0b, \-vmo20\ => \-vmo20\, \-mapi12b\ => \-mapi12b\, \-mapi11b\ => \-mapi11b\, \-mapi10b\ => \-mapi10b\, \-mapi9b\ => \-mapi9b\, \-mapi8b\ => \-mapi8b\, \-vm1wpb\ => \-vm1wpb\, \-vma20\ => \-vma20\, \-vmo21\ => \-vmo21\, \-vma21\ => \-vma21\, \-vmo22\ => \-vmo22\, \-vma22\ => \-vma22\, \-vmo23\ => \-vmo23\, \-vma23\ => \-vma23\, \-vmo16\ => \-vmo16\, \-vma16\ => \-vma16\, \-vmo17\ => \-vmo17\, \-vma17\ => \-vma17\, \-vmo18\ => \-vmo18\, \-vma18\ => \-vma18\, \-vmo19\ => \-vmo19\, \-vma19\ => \-vma19\, \-vmo12\ => \-vmo12\, \-vma12\ => \-vma12\, \-vmo13\ => \-vmo13\, \-vma13\ => \-vma13\, \-vmo14\ => \-vmo14\, \-vma14\ => \-vma14\, \-vmo15\ => \-vmo15\, \-vma15\ => \-vma15\, vmoparm => vmoparm, vmopar => vmopar, vm1pari => vm1pari, \-vmap4\ => \-vmap4\, \-vmap3\ => \-vmap3\, \-vmap2\ => \-vmap2\, \-vmap1\ => \-vmap1\, \-vmap0\ => \-vmap0\, \-vmo5\ => \-vmo5\, \-vmo6\ => \-vmo6\, \-vmo7\ => \-vmo7\, \-vmo8\ => \-vmo8\, \-vmo9\ => \-vmo9\, \-vmo10\ => \-vmo10\, \-vmo11\ => \-vmo11\, vmoparl => vmoparl, \-vmo0\ => \-vmo0\, \-vmo1\ => \-vmo1\, \-vmo2\ => \-vmo2\, \-vmo3\ => \-vmo3\, \-vmo4\ => \-vmo4\, vmoparck => vmoparck, vmoparodd => vmoparodd);
  i_vmemdr : entity cadr_book.vmemdr(ttl) port map(\-mapdrive\ => \-mapdrive\, \-pfw\ => \-pfw\, mf24 => mf24, \-pfr\ => \-pfr\, mf25 => mf25, hi12 => hi12, mf26 => mf26, \-vmap4\ => \-vmap4\, mf27 => mf27, \-vmap3\ => \-vmap3\, mf28 => mf28, \-vmap2\ => \-vmap2\, mf29 => mf29, \-vmap1\ => \-vmap1\, mf30 => mf30, \-vmap0\ => \-vmap0\, mf31 => mf31, \-vmo15\ => \-vmo15\, mf8 => mf8, \-vmo14\ => \-vmo14\, mf9 => mf9, \-vmo13\ => \-vmo13\, mf10 => mf10, \-vmo12\ => \-vmo12\, mf11 => mf11, \-vmo11\ => \-vmo11\, mf12 => mf12, \-vmo10\ => \-vmo10\, mf13 => mf13, \-vmo9\ => \-vmo9\, mf14 => mf14, \-vmo8\ => \-vmo8\, mf15 => mf15, \-vmo23\ => \-vmo23\, mf16 => mf16, \-vmo22\ => \-vmo22\, mf17 => mf17, \-vmo21\ => \-vmo21\, mf18 => mf18, \-vmo20\ => \-vmo20\, mf19 => mf19, \-vmo19\ => \-vmo19\, mf20 => mf20, \-vmo18\ => \-vmo18\, mf21 => mf21, \-vmo17\ => \-vmo17\, mf22 => mf22, \-vmo16\ => \-vmo16\, mf23 => mf23, tse1a => tse1a, srcmap => srcmap, \-vmo7\ => \-vmo7\, mf0 => mf0, \-vmo6\ => \-vmo6\, mf1 => mf1, \-vmo5\ => \-vmo5\, mf2 => mf2, \-vmo4\ => \-vmo4\, mf3 => mf3, \-vmo3\ => \-vmo3\, mf4 => mf4, \-vmo2\ => \-vmo2\, mf5 => mf5, \-vmo1\ => \-vmo1\, mf6 => mf6, \-vmo0\ => \-vmo0\, mf7 => mf7, gnd => gnd, \-lvmo23\ => \-lvmo23\, \-lvmo22\ => \-lvmo22\, \-pma21\ => \-pma21\, \-pma20\ => \-pma20\, memstart => memstart, \-pma19\ => \-pma19\, \-pma18\ => \-pma18\, \-pma17\ => \-pma17\, \-pma16\ => \-pma16\, \-pma15\ => \-pma15\, \-pma14\ => \-pma14\, \-pma13\ => \-pma13\, \-pma12\ => \-pma12\, \-pma11\ => \-pma11\, \-pma10\ => \-pma10\, \-pma9\ => \-pma9\, \-pma8\ => \-pma8\, \-vma6\ => \-vma6\, \-vma5\ => \-vma5\, \-vma4\ => \-vma4\, \-vma3\ => \-vma3\, \-vma2\ => \-vma2\, \-vma1\ => \-vma1\, \-vma0\ => \-vma0\, \-vma7\ => \-vma7\, \-adrpar\ => \-adrpar\, \-srcmap\ => \-srcmap\);


--- Memory Control Logic (vctl)
  i_vctl1 : entity cadr_book.vctl1(ttl) port map(\-reset\ => \-reset\, rdcyc => rdcyc, wrcyc => wrcyc, clk2a => clk2a, wmap => wmap, \-wmapd\ => \-wmapd\, wmapd => wmapd, memprepare => memprepare, \-memwr\ => \-memwr\, \-memprepare\ => \-memprepare\, \-lvmo22\ => \-lvmo22\, \-pfw\ => \-pfw\, \-pfr\ => \-pfr\, \-vmaok\ => \-vmaok\, \-mfinishd\ => \-mfinishd\, memrq => memrq, mclk1a => mclk1a, hi11 => hi11, mbusy => mbusy, \rd.in.progress\ => \rd.in.progress\, \set.rd.in.progress\ => \set.rd.in.progress\, \-rdfinish\ => \-rdfinish\, \-mfinish\ => \-mfinish\, clk2c => clk2c, \-memop\ => \-memop\, \-memack\ => \-memack\, \-memrd\ => \-memrd\, \-ifetch\ => \-ifetch\, memstart => memstart, \-memstart\ => \-memstart\, \-mbusy.sync\ => \-mbusy.sync\, \mbusy.sync\ => \mbusy.sync\, hi4 => hi4, destmem => destmem, \-memgrant\ => \-memgrant\, \use.md\ => \use.md\, \-wait\ => \-wait\, gnd => gnd, needfetch => needfetch, lcinc => lcinc, \-hang\ => \-hang\, \-clk3g\ => \-clk3g\);
  i_vctl2 : entity cadr_book.vctl2(ttl) port map(mapwr0d => mapwr0d, \-wmapd\ => \-wmapd\, \-vma26\ => \-vma26\, mapwr1d => mapwr1d, \-vma25\ => \-vma25\, wp1a => wp1a, \-vm0wpa\ => \-vm0wpa\, \-vm0wpb\ => \-vm0wpb\, \-vm1wpa\ => \-vm1wpa\, wp1b => wp1b, \-vm1wpb\ => \-vm1wpb\, \-lvmo23\ => \-lvmo23\, \-pfr\ => \-pfr\, \-wmap\ => \-wmap\, wmap => wmap, \-memrq\ => \-memrq\, memrq => memrq, \-memprepare\ => \-memprepare\, memprepare => memprepare, destmem => destmem, \-destmem\ => \-destmem\, mdsela => mdsela, \-destmdr\ => \-destmdr\, clk2c => clk2c, mdselb => mdselb, \-destvma\ => \-destvma\, \-ifetch\ => \-ifetch\, \-vmaenb\ => \-vmaenb\, hi11 => hi11, vmasela => vmasela, vmaselb => vmaselb, wrcyc => wrcyc, \lm_drive_enb\ => \lm_drive_enb\, \-memdrive.a\ => \-memdrive.a\, \-memdrive.b\ => \-memdrive.b\, \-memwr\ => \-memwr\, \-memrd\ => \-memrd\, ir20 => ir20, ir19 => ir19, \use.md\ => \use.md\, \-srcmd\ => \-srcmd\, nopa => nopa, \-nopa\ => \-nopa\);
  i_olord1 : entity icmem_book.olord1(ttl) port map(\-clock_reset_a\ => \-clock_reset_a\, speed1a => speed1a, sspeed1 => sspeed1, speedclk => speedclk, sspeed0 => sspeed0, speed0a => speed0a, speed1 => speed1, speed0 => speed0, \-reset\ => \-reset\, spy0 => spy0, spy1 => spy1, spy2 => spy2, errstop => errstop, \-ldmode\ => \-ldmode\, stathenb => stathenb, spy3 => spy3, trapenb => trapenb, spy4 => spy4, spy5 => spy5, promdisable => promdisable, \-opcinh\ => \-opcinh\, opcinh => opcinh, \-ldopc\ => \-ldopc\, opcclk => opcclk, \-opcclk\ => \-opcclk\, \-lpc.hold\ => \-lpc.hold\, \lpc.hold\ => \lpc.hold\, ldstat => ldstat, \-ldstat\ => \-ldstat\, \-idebug\ => \-idebug\, idebug => idebug, \-ldclk\ => \-ldclk\, nop11 => nop11, \-nop11\ => \-nop11\, \-step\ => \-step\, step => step, promdisabled => promdisabled, sstep => sstep, ssdone => ssdone, mclk5a => mclk5a, srun => srun, run => run, \-boot\ => \-boot\, \-run\ => \-run\, \-ssdone\ => \-ssdone\, \-errhalt\ => \-errhalt\, \-wait\ => \-wait\, \-stathalt\ => \-stathalt\, machrun => machrun, \stat.ovf\ => \stat.ovf\, \-stc32\ => \-stc32\, \-tpr60\ => \-tpr60\, gnd => gnd, statstop => statstop, \-machruna\ => \-machruna\, \-machrun\ => \-machrun\);
  i_olord2 : entity icmem_book.olord2(ttl) port map(\-ape\ => \-ape\, \-mpe\ => \-mpe\, \-pdlpe\ => \-pdlpe\, \-dpe\ => \-dpe\, \-ipe\ => \-ipe\, \-spe\ => \-spe\, \-higherr\ => \-higherr\, err => err, \-mempe\ => \-mempe\, \-v0pe\ => \-v0pe\, \-v1pe\ => \-v1pe\, \-halted\ => \-halted\, hi1 => hi1, gnd => gnd, aparok => aparok, mmemparok => mmemparok, pdlparok => pdlparok, dparok => dparok, clk5a => clk5a, iparok => iparok, spcparok => spcparok, highok => highok, memparok => memparok, v0parok => v0parok, vmoparok => vmoparok, statstop => statstop, \stat.ovf\ => \stat.ovf\, \-halt\ => \-halt\, \-mclk5\ => \-mclk5\, mclk5a => mclk5a, \-clk5\ => \-clk5\, \-reset\ => \-reset\, reset => reset, \bus.power.reset_l\ => \bus.power.reset_l\, \power_reset_a\ => \power_reset_a\, \-upperhighok\ => \-upperhighok\, \-lowerhighok\ => \-lowerhighok\, \-boot\ => \-boot\, \prog.bus.reset\ => \prog.bus.reset\, \-bus.reset\ => \-bus.reset\, \-clock_reset_b\ => \-clock_reset_b\, \-clock_reset_a\ => \-clock_reset_a\, \-power_reset\ => \-power_reset\, srun => srun, \boot.trap\ => \boot.trap\, hi2 => hi2, \-boot1\ => \-boot1\, \-boot2\ => \-boot2\, \-ldmode\ => \-ldmode\, ldmode => ldmode, mclk5 => mclk5, clk5 => clk5, \-busint.lm.reset\ => \-busint.lm.reset\, \-prog.reset\ => \-prog.reset\, spy6 => spy6, \-errhalt\ => \-errhalt\, errstop => errstop, \prog.boot\ => \prog.boot\, spy7 => spy7);


--- Other (...)
  i_stat : entity icmem_book.stat(ttl) port map(hi1 => hi1, clk5a => clk5a, iwr12 => iwr12, iwr13 => iwr13, iwr14 => iwr14, iwr15 => iwr15, gnd => gnd, \-ldstat\ => \-ldstat\, \-stc12\ => \-stc12\, st15 => st15, st14 => st14, st13 => st13, st12 => st12, \-stc16\ => \-stc16\, iwr16 => iwr16, iwr17 => iwr17, iwr18 => iwr18, iwr19 => iwr19, st19 => st19, st18 => st18, st17 => st17, st16 => st16, \-stc20\ => \-stc20\, iwr20 => iwr20, iwr21 => iwr21, iwr22 => iwr22, iwr23 => iwr23, st23 => st23, st22 => st22, st21 => st21, st20 => st20, \-stc24\ => \-stc24\, iwr24 => iwr24, iwr25 => iwr25, iwr26 => iwr26, iwr27 => iwr27, st27 => st27, st26 => st26, st25 => st25, st24 => st24, \-stc28\ => \-stc28\, iwr28 => iwr28, iwr29 => iwr29, iwr30 => iwr30, iwr31 => iwr31, st31 => st31, st30 => st30, st29 => st29, st28 => st28, \-stc32\ => \-stc32\, \-spy.sth\ => \-spy.sth\, spy8 => spy8, spy9 => spy9, spy10 => spy10, spy11 => spy11, spy12 => spy12, spy13 => spy13, spy14 => spy14, spy15 => spy15, spy0 => spy0, spy1 => spy1, spy2 => spy2, spy3 => spy3, spy4 => spy4, spy5 => spy5, spy6 => spy6, spy7 => spy7, \-spy.stl\ => \-spy.stl\, st11 => st11, st10 => st10, st9 => st9, st8 => st8, st7 => st7, st6 => st6, st5 => st5, st4 => st4, st3 => st3, st2 => st2, st1 => st1, st0 => st0, iwr0 => iwr0, iwr1 => iwr1, iwr2 => iwr2, iwr3 => iwr3, \-statbit\ => \-statbit\, \-stc4\ => \-stc4\, iwr4 => iwr4, iwr5 => iwr5, iwr6 => iwr6, iwr7 => iwr7, \-stc8\ => \-stc8\, iwr8 => iwr8, iwr9 => iwr9, iwr10 => iwr10, iwr11 => iwr11);
  i_opcs : entity icmem_book.opcs(ttl) port map(hi2 => hi2, opc13 => opc13, gnd => gnd, pc13 => pc13, opcinha => opcinha, opcclka => opcclka, pc12 => pc12, opc12 => opc12, opc11 => opc11, pc11 => pc11, pc10 => pc10, opc10 => opc10, opc9 => opc9, pc9 => pc9, opcclkc => opcclkc, pc8 => pc8, opc8 => opc8, opc7 => opc7, pc7 => pc7, pc6 => pc6, opc6 => opc6, \-opcinh\ => \-opcinh\, opcinhb => opcinhb, opc5 => opc5, pc5 => pc5, opcclkb => opcclkb, pc4 => pc4, opc4 => opc4, opc3 => opc3, pc3 => pc3, pc2 => pc2, opc2 => opc2, opc1 => opc1, pc1 => pc1, pc0 => pc0, opc0 => opc0, \-clk5\ => \-clk5\, opcclk => opcclk);
  i_iwrpar : entity icmem_book.iwrpar(ttl) port map(iwr41 => iwr41, iwr42 => iwr42, iwr43 => iwr43, iwr44 => iwr44, iwr45 => iwr45, iwr46 => iwr46, iwr47 => iwr47, iwrp4 => iwrp4, iwr36 => iwr36, iwr37 => iwr37, iwr38 => iwr38, iwr39 => iwr39, iwr40 => iwr40, iwr29 => iwr29, iwr30 => iwr30, iwr31 => iwr31, iwr32 => iwr32, iwr33 => iwr33, iwr34 => iwr34, iwr35 => iwr35, iwrp3 => iwrp3, iwr24 => iwr24, iwr25 => iwr25, iwr26 => iwr26, iwr27 => iwr27, iwr28 => iwr28, iwr17 => iwr17, iwr18 => iwr18, iwr19 => iwr19, iwr20 => iwr20, iwr21 => iwr21, iwr22 => iwr22, iwr23 => iwr23, iwrp2 => iwrp2, iwr12 => iwr12, iwr13 => iwr13, iwr14 => iwr14, iwr15 => iwr15, iwr16 => iwr16, iwr5 => iwr5, iwr6 => iwr6, iwr7 => iwr7, iwr8 => iwr8, iwr9 => iwr9, iwr10 => iwr10, iwr11 => iwr11, iwrp1 => iwrp1, iwr0 => iwr0, iwr1 => iwr1, iwr2 => iwr2, iwr3 => iwr3, iwr4 => iwr4, gnd => gnd, iwr48 => iwr48);
  i_trap : entity cadr_book.trap(ttl) port map(mdparerr => mdparerr, mdpareven => mdpareven, mdpar => mdpar, \-md5\ => \-md5\, \-md6\ => \-md6\, \-md7\ => \-md7\, \-md8\ => \-md8\, \-md9\ => \-md9\, \-md10\ => \-md10\, \-md11\ => \-md11\, mdparl => mdparl, \-md0\ => \-md0\, \-md1\ => \-md1\, \-md2\ => \-md2\, \-md3\ => \-md3\, \-md4\ => \-md4\, \-md17\ => \-md17\, \-md18\ => \-md18\, \-md19\ => \-md19\, \-md20\ => \-md20\, \-md21\ => \-md21\, \-md22\ => \-md22\, \-md23\ => \-md23\, mdparm => mdparm, \-md12\ => \-md12\, \-md13\ => \-md13\, \-md14\ => \-md14\, \-md15\ => \-md15\, \-md16\ => \-md16\, \-md29\ => \-md29\, \-md30\ => \-md30\, \-md31\ => \-md31\, gnd => gnd, mdparodd => mdparodd, \-md24\ => \-md24\, \-md25\ => \-md25\, \-md26\ => \-md26\, \-md27\ => \-md27\, \-md28\ => \-md28\, mdhaspar => mdhaspar, \use.md\ => \use.md\, \-wait\ => \-wait\, \-parerr\ => \-parerr\, \-trap\ => \-trap\, \boot.trap\ => \boot.trap\, \-trapenb\ => \-trapenb\, trapenb => trapenb, \-memparok\ => \-memparok\, trapb => trapb, trapa => trapa, memparok => memparok);
  i_spy0 : entity icmem_book.spy0(ttl) port map(eadr0 => eadr0, eadr1 => eadr1, eadr2 => eadr2, \-dbread\ => \-dbread\, eadr3 => eadr3, hi1 => hi1, \-spy.obh\ => \-spy.obh\, \-spy.obl\ => \-spy.obl\, \-spy.pc\ => \-spy.pc\, \-spy.opc\ => \-spy.opc\, \-spy.irh\ => \-spy.irh\, \-spy.irm\ => \-spy.irm\, \-spy.irl\ => \-spy.irl\, gnd => gnd, \-spy.sth\ => \-spy.sth\, \-spy.stl\ => \-spy.stl\, \-spy.ah\ => \-spy.ah\, \-spy.al\ => \-spy.al\, \-spy.mh\ => \-spy.mh\, \-spy.ml\ => \-spy.ml\, \-spy.flag2\ => \-spy.flag2\, \-spy.flag1\ => \-spy.flag1\, \-dbwrite\ => \-dbwrite\, \-ldmode\ => \-ldmode\, \-ldopc\ => \-ldopc\, \-ldclk\ => \-ldclk\, \-lddbirh\ => \-lddbirh\, \-lddbirm\ => \-lddbirm\, \-lddbirl\ => \-lddbirl\);
  i_spy1 : entity cadr_book.spy1(ttl) port map(\-spy.obl\ => \-spy.obl\, ob7 => ob7, spy0 => spy0, ob6 => ob6, spy1 => spy1, ob5 => ob5, spy2 => spy2, ob4 => ob4, spy3 => spy3, ob3 => ob3, spy4 => spy4, ob2 => ob2, spy5 => spy5, ob1 => ob1, spy6 => spy6, ob0 => ob0, spy7 => spy7, ob15 => ob15, spy8 => spy8, ob14 => ob14, spy9 => spy9, ob13 => ob13, spy10 => spy10, ob12 => ob12, spy11 => spy11, ob11 => ob11, spy12 => spy12, ob10 => ob10, spy13 => spy13, ob9 => ob9, spy14 => spy14, ob8 => ob8, spy15 => spy15, \-spy.obh\ => \-spy.obh\, ob23 => ob23, ob22 => ob22, ob21 => ob21, ob20 => ob20, ob19 => ob19, ob18 => ob18, ob17 => ob17, ob16 => ob16, ob31 => ob31, ob30 => ob30, ob29 => ob29, ob28 => ob28, ob27 => ob27, ob26 => ob26, ob25 => ob25, ob24 => ob24, \-spy.irl\ => \-spy.irl\, ir7 => ir7, ir6 => ir6, ir5 => ir5, ir4 => ir4, ir3 => ir3, ir2 => ir2, ir1 => ir1, ir0 => ir0, ir15 => ir15, ir14 => ir14, ir13 => ir13, ir12 => ir12, ir11 => ir11, ir10 => ir10, ir9 => ir9, ir8 => ir8, \-spy.irh\ => \-spy.irh\, ir47 => ir47, ir46 => ir46, ir45 => ir45, ir44 => ir44, ir43 => ir43, ir42 => ir42, ir41 => ir41, ir40 => ir40, ir39 => ir39, ir38 => ir38, ir37 => ir37, ir36 => ir36, ir35 => ir35, ir34 => ir34, ir33 => ir33, ir32 => ir32, \-spy.irm\ => \-spy.irm\, ir31 => ir31, ir30 => ir30, ir29 => ir29, ir28 => ir28, ir27 => ir27, ir26 => ir26, ir25 => ir25, ir24 => ir24, ir23 => ir23, ir22 => ir22, ir21 => ir21, ir20 => ir20, ir19 => ir19, ir18 => ir18, ir17 => ir17, ir16 => ir16);
  i_spy2 : entity cadr_book.spy2(ttl) port map(\-spy.al\ => \-spy.al\, aa15 => aa15, spy8 => spy8, aa14 => aa14, spy9 => spy9, aa13 => aa13, spy10 => spy10, aa12 => aa12, spy11 => spy11, aa11 => aa11, spy12 => spy12, aa10 => aa10, spy13 => spy13, aa9 => aa9, spy14 => spy14, aa8 => aa8, spy15 => spy15, aa7 => aa7, spy0 => spy0, aa6 => aa6, spy1 => spy1, aa5 => aa5, spy2 => spy2, aa4 => aa4, spy3 => spy3, aa3 => aa3, spy4 => spy4, aa2 => aa2, spy5 => spy5, aa1 => aa1, spy6 => spy6, aa0 => aa0, spy7 => spy7, \-spy.ah\ => \-spy.ah\, a31a => a31a, a30 => a30, a29 => a29, a28 => a28, a27 => a27, a26 => a26, a25 => a25, a24 => a24, a23 => a23, a22 => a22, a21 => a21, a20 => a20, a19 => a19, a18 => a18, a17 => a17, a16 => a16, \-spy.flag2\ => \-spy.flag2\, ir48 => ir48, nop => nop, \-vmaok\ => \-vmaok\, jcond => jcond, pcs1 => pcs1, pcs0 => pcs0, wmapd => wmapd, destspcd => destspcd, iwrited => iwrited, imodd => imodd, pdlwrited => pdlwrited, spushd => spushd, \-spy.ml\ => \-spy.ml\, m15 => m15, m14 => m14, m13 => m13, m12 => m12, m11 => m11, m10 => m10, m9 => m9, m8 => m8, m7 => m7, m6 => m6, m5 => m5, m4 => m4, m3 => m3, m2 => m2, m1 => m1, m0 => m0, \-spy.mh\ => \-spy.mh\, m23 => m23, m22 => m22, m21 => m21, m20 => m20, m19 => m19, m18 => m18, m17 => m17, m16 => m16, m31 => m31, m30 => m30, m29 => m29, m28 => m28, m27 => m27, m26 => m26, m25 => m25, m24 => m24);
  i_spy4 : entity icmem_book.spy4(ttl) port map(\-spy.flag1\ => \-spy.flag1\, \-wait\ => \-wait\, spy8 => spy8, \-v1pe\ => \-v1pe\, spy9 => spy9, \-v0pe\ => \-v0pe\, spy10 => spy10, promdisable => promdisable, spy11 => spy11, \-stathalt\ => \-stathalt\, spy12 => spy12, err => err, spy13 => spy13, ssdone => ssdone, spy14 => spy14, srun => srun, spy15 => spy15, \-higherr\ => \-higherr\, spy0 => spy0, \-mempe\ => \-mempe\, spy1 => spy1, \-ipe\ => \-ipe\, spy2 => spy2, \-dpe\ => \-dpe\, spy3 => spy3, \-spe\ => \-spe\, spy4 => spy4, \-pdlpe\ => \-pdlpe\, spy5 => spy5, \-mpe\ => \-mpe\, spy6 => spy6, \-ape\ => \-ape\, spy7 => spy7, \-spy.pc\ => \-spy.pc\, gnd => gnd, pc13 => pc13, pc12 => pc12, pc11 => pc11, pc10 => pc10, pc9 => pc9, pc8 => pc8, pc7 => pc7, pc6 => pc6, pc5 => pc5, pc4 => pc4, pc3 => pc3, pc2 => pc2, pc1 => pc1, pc0 => pc0, \-spy.opc\ => \-spy.opc\, opc13 => opc13, opc12 => opc12, opc11 => opc11, opc10 => opc10, opc9 => opc9, opc8 => opc8, opc7 => opc7, opc6 => opc6, opc5 => opc5, opc4 => opc4, opc3 => opc3, opc2 => opc2, opc1 => opc1, opc0 => opc0);
  i_opcd : entity cadr_book.opcd(ttl) port map(\-srcdc\ => \-srcdc\, \-srcopc\ => \-srcopc\, \-opcdrive\ => \-opcdrive\, opc7 => opc7, mf4 => mf4, opc6 => opc6, mf5 => mf5, opc5 => opc5, mf6 => mf6, opc4 => opc4, mf7 => mf7, dc7 => dc7, dc6 => dc6, dc5 => dc5, dc4 => dc4, dcdrive => dcdrive, opc3 => opc3, mf0 => mf0, opc2 => opc2, mf1 => mf1, opc1 => opc1, mf2 => mf2, opc0 => opc0, mf3 => mf3, dc3 => dc3, dc2 => dc2, dc1 => dc1, dc0 => dc0, tse1b => tse1b, \-zero16.drive\ => \-zero16.drive\, zero16 => zero16, \zero16.drive\ => \zero16.drive\, \zero12.drive\ => \zero12.drive\, gnd => gnd, mf24 => mf24, mf25 => mf25, mf26 => mf26, mf27 => mf27, mf28 => mf28, mf29 => mf29, mf30 => mf30, mf31 => mf31, mf16 => mf16, mf17 => mf17, mf18 => mf18, mf19 => mf19, mf20 => mf20, mf21 => mf21, mf22 => mf22, mf23 => mf23, mf12 => mf12, mf13 => mf13, opc13 => opc13, mf14 => mf14, opc12 => opc12, mf15 => mf15, opc11 => opc11, mf8 => mf8, opc10 => opc10, mf9 => mf9, opc9 => opc9, mf10 => mf10, opc8 => opc8, mf11 => mf11, dc9 => dc9, dc8 => dc8, \-srcpdlidx\ => \-srcpdlidx\, \-srcpdlptr\ => \-srcpdlptr\);
  i_mo0 : entity cadr_book.mo0(ttl) port map(alu15 => alu15, r15 => r15, a15 => a15, ob15 => ob15, gnd => gnd, osel1b => osel1b, osel0b => osel0b, msk15 => msk15, alu14 => alu14, alu16 => alu16, r14 => r14, a14 => a14, ob14 => ob14, msk14 => msk14, alu13 => alu13, r13 => r13, a13 => a13, ob13 => ob13, msk13 => msk13, alu12 => alu12, r12 => r12, a12 => a12, ob12 => ob12, msk12 => msk12, alu11 => alu11, alu7 => alu7, r7 => r7, a7 => a7, ob7 => ob7, msk7 => msk7, alu6 => alu6, alu8 => alu8, r6 => r6, a6 => a6, ob6 => ob6, msk6 => msk6, alu5 => alu5, r5 => r5, a5 => a5, ob5 => ob5, msk5 => msk5, alu4 => alu4, r4 => r4, a4 => a4, ob4 => ob4, msk4 => msk4, alu3 => alu3, r11 => r11, a11 => a11, ob11 => ob11, msk11 => msk11, alu10 => alu10, r10 => r10, a10 => a10, ob10 => ob10, msk10 => msk10, alu9 => alu9, r3 => r3, a3 => a3, ob3 => ob3, msk3 => msk3, alu2 => alu2, r2 => r2, a2 => a2, ob2 => ob2, msk2 => msk2, alu1 => alu1, r9 => r9, a9 => a9, ob9 => ob9, msk9 => msk9, r8 => r8, a8 => a8, ob8 => ob8, msk8 => msk8, r1 => r1, a1 => a1, ob1 => ob1, msk1 => msk1, alu0 => alu0, r0 => r0, a0 => a0, ob0 => ob0, msk0 => msk0, q31 => q31);
  i_mo1 : entity cadr_book.mo1(ttl) port map(alu31 => alu31, r31 => r31, a31b => a31b, ob31 => ob31, gnd => gnd, osel1a => osel1a, osel0a => osel0a, msk31 => msk31, alu30 => alu30, alu32 => alu32, r30 => r30, a30 => a30, ob30 => ob30, msk30 => msk30, alu29 => alu29, r29 => r29, a29 => a29, ob29 => ob29, msk29 => msk29, alu28 => alu28, r28 => r28, a28 => a28, ob28 => ob28, msk28 => msk28, alu27 => alu27, alu23 => alu23, r23 => r23, a23 => a23, ob23 => ob23, msk23 => msk23, alu22 => alu22, alu24 => alu24, r22 => r22, a22 => a22, ob22 => ob22, msk22 => msk22, alu21 => alu21, r21 => r21, a21 => a21, ob21 => ob21, msk21 => msk21, alu20 => alu20, r20 => r20, a20 => a20, ob20 => ob20, msk20 => msk20, alu19 => alu19, r27 => r27, a27 => a27, ob27 => ob27, msk27 => msk27, alu26 => alu26, r24 => r24, a24 => a24, ob24 => ob24, msk24 => msk24, alu25 => alu25, r26 => r26, a26 => a26, ob26 => ob26, msk26 => msk26, r25 => r25, a25 => a25, ob25 => ob25, msk25 => msk25, r19 => r19, a19 => a19, ob19 => ob19, msk19 => msk19, alu18 => alu18, r18 => r18, a18 => a18, ob18 => ob18, msk18 => msk18, alu17 => alu17, r17 => r17, a17 => a17, ob17 => ob17, msk17 => msk17, alu16 => alu16, r16 => r16, a16 => a16, ob16 => ob16, msk16 => msk16, alu15 => alu15);
  i_bcterm : entity cadr_book.bcterm(ttl) port map(mem0 => mem0, mem1 => mem1, mem2 => mem2, mem3 => mem3, mem4 => mem4, mem5 => mem5, mem12 => mem12, mem13 => mem13, mem14 => mem14, mem15 => mem15, mem16 => mem16, mem17 => mem17, mem24 => mem24, mem25 => mem25, mem26 => mem26, mem27 => mem27, mem28 => mem28, mem29 => mem29, \-memgrant\ => \-memgrant\, int => int, \-loadmd\ => \-loadmd\, \-ignpar\ => \-ignpar\, \-memack\ => \-memack\);
  i_ipar : entity cadr_book.ipar(ttl) port map(ir41 => ir41, ir42 => ir42, ir43 => ir43, ir44 => ir44, ir45 => ir45, ir46 => ir46, ir47 => ir47, ipar3 => ipar3, ir36 => ir36, ir37 => ir37, ir38 => ir38, ir39 => ir39, ir40 => ir40, ir5 => ir5, ir6 => ir6, ir7 => ir7, ir8 => ir8, ir9 => ir9, ir10 => ir10, ir11 => ir11, ipar0 => ipar0, ir0 => ir0, ir1 => ir1, ir2 => ir2, ir3 => ir3, ir4 => ir4, ir29 => ir29, ir30 => ir30, ir31 => ir31, ir32 => ir32, ir33 => ir33, ir34 => ir34, ir35 => ir35, ipar2 => ipar2, ir24 => ir24, ir25 => ir25, ir26 => ir26, ir27 => ir27, ir28 => ir28, gnd => gnd, iparity => iparity, ipar1 => ipar1, ir48 => ir48, ir17 => ir17, ir18 => ir18, ir19 => ir19, ir20 => ir20, ir21 => ir21, ir22 => ir22, ir23 => ir23, ir12 => ir12, ir13 => ir13, ir14 => ir14, ir15 => ir15, ir16 => ir16, imodd => imodd, iparok => iparok);

  gnd <= '0';

  -- Manual Overlord.

  speed0   <= '0';
  speed1   <= '0';
  \-ilong\ <= not '0';
  
  process
  begin
    \-hang\          <= not '0';
    \-clock_reset_b\ <= not '0';
    wait for 20 ns;
    \-clock_reset_b\ <= not '1';
    wait;
  end process;
  
  -- Poor substitute for the 5 octal display that was on the lower
  -- left-hand corner of the front door on the CADR.  See the PCTL
  -- prints.
  process (cyclecompleted)
    variable cycles : integer := 0;
  begin
    if rising_edge(cyclecompleted) then
      cycles := cycles + 1;
      
--      report integer'image(cycles) & ": PC:" & to_hstring(pc);
      if tilt1 then report "TILT1"; end if;
      if tilt0 then report "TILT0"; end if;
      if dpe then report "DPE"; end if;
      if ipe then report "IPE"; end if;
      if promenable then report "PROMENABLE"; end if;
    end if;
    
    if cycles >= 1000 then
      finish;
    end if;
  end process;
  
end architecture;
