-- CADR1_BUSPAR
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_buspar is
  port (
    \bus 0\ : in std_logic;
    \bus 0-11 par odd\ : inout std_logic;
    \bus 1\ : in std_logic;
    \bus 10\ : in std_logic;
    \bus 11\ : in std_logic;
    \bus 12\ : in std_logic;
    \bus 12-23 par odd\ : inout std_logic;
    \bus 13\ : in std_logic;
    \bus 14\ : in std_logic;
    \bus 15\ : in std_logic;
    \bus 16\ : in std_logic;
    \bus 17\ : in std_logic;
    \bus 18\ : in std_logic;
    \bus 19\ : in std_logic;
    \bus 2\ : in std_logic;
    \bus 20\ : in std_logic;
    \bus 21\ : in std_logic;
    \bus 22\ : in std_logic;
    \bus 23\ : in std_logic;
    \bus 24\ : in std_logic;
    \bus 25\ : in std_logic;
    \bus 26\ : in std_logic;
    \bus 27\ : in std_logic;
    \bus 28\ : in std_logic;
    \bus 29\ : in std_logic;
    \bus 3\ : in std_logic;
    \bus 30\ : in std_logic;
    \bus 31\ : in std_logic;
    \bus 4\ : in std_logic;
    \bus 5\ : in std_logic;
    \bus 6\ : in std_logic;
    \bus 7\ : in std_logic;
    \bus 8\ : in std_logic;
    \bus 9\ : in std_logic;
    \bus par even\ : out std_logic;
    \bus par odd\ : out std_logic
  );
end entity;
