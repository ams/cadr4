-- IRAM21 -- RAM 4K-8K, 24-35

library work;
use work.dip.all;
use work.misc.all;

architecture behv of cadr_iram21 is
begin
iram21_1a26 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i31, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr31, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1a27 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i32, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr32, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1a28 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i33, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr33, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1a29 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i34, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr34, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1a30 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i35, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr35, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1b26 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i26, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr26, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1b27 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i27, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr27, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1b28 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i28, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr28, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1b29 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i29, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr29, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1b30 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i30, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr30, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1c27 : dip_74s04a port map (p1 => \-pcc6\, p2 => pc6j, p3 => \-pcc7\, p4 => pc7j, p5 => \-pcc8\, p6 => pc8j, p8 => pc9j, p9 => \-pcc9\, p10 => pc10j, p11 => \-pcc10\, p12 => pc11j, p13 => \-pcc11\);
iram21_1c28 : dip_74s04a port map (p1 => \-pcc0\, p2 => pc0j, p3 => \-pcc1\, p4 => pc1j, p5 => \-pcc2\, p6 => pc2j, p8 => pc3j, p9 => \-pcc3\, p10 => pc4j, p11 => \-pcc4\, p12 => pc5j, p13 => \-pcc5\);
iram21_1c29 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i24, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr24, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
iram21_1c30 : dip_2147 port map (p1 => pc0j, p2 => pc1j, p3 => pc2j, p4 => pc3j, p5 => pc4j, p6 => pc5j, p7 => i25, p8 => \-iwej\, p10 => \-ice1c\, p11 => iwr25, p12 => pc11j, p13 => pc10j, p14 => pc9j, p15 => pc8j, p16 => pc7j, p17 => pc6j);
end architecture;
