-- CADR1_WBUF
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_wbuf is
  port (
    \-ubpn0a\ : inout std_logic;
    \-ubpn0b\ : inout std_logic;
    \-ubpn1a\ : inout std_logic;
    \-ubpn1b\ : inout std_logic;
    \-ubpn2a\ : inout std_logic;
    \-ubpn2b\ : inout std_logic;
    \-ubpn3a\ : inout std_logic;
    \-ubpn3b\ : inout std_logic;
    \-wbufwe\ : inout std_logic;
    udi0 : inout std_logic;
    udi1 : inout std_logic;
    udi10 : inout std_logic;
    udi11 : inout std_logic;
    udi12 : inout std_logic;
    udi13 : inout std_logic;
    udi14 : inout std_logic;
    udi15 : inout std_logic;
    udi2 : inout std_logic;
    udi3 : inout std_logic;
    udi4 : inout std_logic;
    udi5 : inout std_logic;
    udi6 : inout std_logic;
    udi7 : inout std_logic;
    udi8 : inout std_logic;
    udi9 : inout std_logic;
    wbuf0 : inout std_logic;
    wbuf1 : inout std_logic;
    wbuf10 : inout std_logic;
    wbuf11 : inout std_logic;
    wbuf12 : inout std_logic;
    wbuf13 : inout std_logic;
    wbuf14 : inout std_logic;
    wbuf15 : inout std_logic;
    wbuf2 : inout std_logic;
    wbuf3 : inout std_logic;
    wbuf4 : inout std_logic;
    wbuf5 : inout std_logic;
    wbuf6 : inout std_logic;
    wbuf7 : inout std_logic;
    wbuf8 : inout std_logic;
    wbuf9 : inout std_logic
  );
end entity;
