library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_16dummy is
  port (
    dummy : in std_logic
    );
end ic_16dummy;

architecture ttl of ic_16dummy is
begin

end ttl;
