library ieee;
use ieee.std_logic_1164.all;

entity apar is
  port (
    a26       : in  std_logic;
    a27       : in  std_logic;
    a28       : in  std_logic;
    a29       : in  std_logic;
    a30       : in  std_logic;
    a31b      : in  std_logic;
    aparity   : in  std_logic;
    aparok    : out std_logic;
    aparl     : out std_logic;
    aparm     : out std_logic;
    gnd       : in  std_logic;
    a24       : in  std_logic;
    a25       : in  std_logic;
    a17       : in  std_logic;
    a18       : in  std_logic;
    a19       : in  std_logic;
    a20       : in  std_logic;
    a21       : in  std_logic;
    a22       : in  std_logic;
    a23       : in  std_logic;
    a12       : in  std_logic;
    a13       : in  std_logic;
    a14       : in  std_logic;
    a15       : in  std_logic;
    a16       : in  std_logic;
    a5        : in  std_logic;
    a6        : in  std_logic;
    a7        : in  std_logic;
    a8        : in  std_logic;
    a9        : in  std_logic;
    a10       : in  std_logic;
    a11       : in  std_logic;
    a0        : in  std_logic;
    a1        : in  std_logic;
    a2        : in  std_logic;
    a3        : in  std_logic;
    a4        : in  std_logic;
    m17       : in  std_logic;
    m18       : in  std_logic;
    m19       : in  std_logic;
    m20       : in  std_logic;
    m21       : in  std_logic;
    m22       : in  std_logic;
    m23       : in  std_logic;
    mparm     : out std_logic;
    m12       : in  std_logic;
    m13       : in  std_logic;
    m14       : in  std_logic;
    m15       : in  std_logic;
    m16       : in  std_logic;
    m5        : in  std_logic;
    m6        : in  std_logic;
    m7        : in  std_logic;
    m8        : in  std_logic;
    m9        : in  std_logic;
    m10       : in  std_logic;
    m11       : in  std_logic;
    mparl     : out std_logic;
    m0        : in  std_logic;
    m1        : in  std_logic;
    m2        : in  std_logic;
    m3        : in  std_logic;
    m4        : in  std_logic;
    mpareven  : out std_logic;
    srcm      : in  std_logic;
    mmemparok : out std_logic;
    pdlenb    : in  std_logic;
    pdlparok  : out std_logic;
    m26       : in  std_logic;
    m27       : in  std_logic;
    m28       : in  std_logic;
    m29       : in  std_logic;
    m30       : in  std_logic;
    m31       : in  std_logic;
    mparity   : in  std_logic;
    mparodd   : out std_logic;
    m24       : in  std_logic;
    m25       : in  std_logic);
end;
