library ieee;
use ieee.std_logic_1164.all;

entity dip_dummy4 is port (
  p2  : out std_logic;                  -- vco cap2
  p3  : out std_logic                   -- vco cap1
  );
end entity;

architecture empty of dip_dummy4 is
begin
end architecture;