library ieee;
use ieee.std_logic_1164.all;

entity dram1 is
  port (
    wp2         : in  std_logic;
    dispwr      : in  std_logic;
    \-dweb\     : out std_logic;
    \-vmo19\    : out std_logic;
    vmo19       : out std_logic;
    \-vmo18\    : out std_logic;
    vmo18       : out std_logic;
    \-dadr9b\   : out std_logic;
    ir21b       : out std_logic;
    \-dadr8b\   : out std_logic;
    ir20b       : out std_logic;
    \-dadr7b\   : out std_logic;
    ir19b       : in  std_logic;
    ir12b       : in  std_logic;
    ir9b        : out std_logic;
    r0          : in  std_logic;
    dmask0      : in  std_logic;
    \-dmapbenb\ : in  std_logic;
    \-dadr0b\   : out std_logic;
    ir8b        : out std_logic;
    hi6         : in  std_logic;
    dadr10a     : in  std_logic;
    \-dadr1b\   : out std_logic;
    \-dadr2b\   : out std_logic;
    \-dadr3b\   : out std_logic;
    \-dadr4b\   : out std_logic;
    dpc11       : out std_logic;
    \-dadr5b\   : out std_logic;
    \-dadr6b\   : out std_logic;
    aa11        : in  std_logic;
    \-dadr10a\  : in  std_logic;
    dpc10       : out std_logic;
    aa10        : in  std_logic;
    r3          : in  std_logic;
    ir18b       : in  std_logic;
    dmask6      : in  std_logic;
    r6          : in  std_logic;
    ir15b       : in  std_logic;
    dmask3      : in  std_logic;
    dpc9        : out std_logic;
    aa9         : in  std_logic;
    dadr10c     : in  std_logic;
    dpc8        : out std_logic;
    aa8         : in  std_logic;
    \-dadr10c\  : in  std_logic;
    r2          : in  std_logic;
    ir17b       : in  std_logic;
    dmask5      : in  std_logic;
    r5          : in  std_logic;
    ir14b       : in  std_logic;
    dmask2      : in  std_logic;
    dpc7        : out std_logic;
    aa7         : in  std_logic;
    dpc6        : out std_logic;
    aa6         : in  std_logic;
    r1          : in  std_logic;
    ir16b       : in  std_logic;
    dmask4      : in  std_logic;
    r4          : in  std_logic;
    ir13b       : in  std_logic;
    dmask1      : in  std_logic;
    gnd         : in  std_logic;
    ir20        : in  std_logic;
    ir21        : in  std_logic;
    ir22        : in  std_logic;
    ir8         : in  std_logic;
    ir9         : in  std_logic;
    ir22b       : out std_logic);
end;
