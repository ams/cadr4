-- CADR1_XD
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_xd is
  port (
    \-xbus ignpar\ : inout std_logic;
    \-xbus par\ : inout std_logic;
    \-xbus wr\ : inout std_logic;
    \-xbus0\ : inout std_logic;
    \-xbus1\ : inout std_logic;
    \-xbus10\ : inout std_logic;
    \-xbus11\ : inout std_logic;
    \-xbus12\ : inout std_logic;
    \-xbus13\ : inout std_logic;
    \-xbus14\ : inout std_logic;
    \-xbus15\ : inout std_logic;
    \-xbus16\ : inout std_logic;
    \-xbus17\ : inout std_logic;
    \-xbus18\ : inout std_logic;
    \-xbus19\ : inout std_logic;
    \-xbus2\ : inout std_logic;
    \-xbus20\ : inout std_logic;
    \-xbus21\ : inout std_logic;
    \-xbus22\ : inout std_logic;
    \-xbus23\ : inout std_logic;
    \-xbus24\ : inout std_logic;
    \-xbus25\ : inout std_logic;
    \-xbus26\ : inout std_logic;
    \-xbus27\ : inout std_logic;
    \-xbus28\ : inout std_logic;
    \-xbus29\ : inout std_logic;
    \-xbus3\ : inout std_logic;
    \-xbus30\ : inout std_logic;
    \-xbus31\ : inout std_logic;
    \-xbus4\ : inout std_logic;
    \-xbus5\ : inout std_logic;
    \-xbus6\ : inout std_logic;
    \-xbus7\ : inout std_logic;
    \-xbus8\ : inout std_logic;
    \-xbus9\ : inout std_logic;
    \-xdrive\ : inout std_logic;
    bus0 : inout std_logic;
    bus1 : inout std_logic;
    bus10 : inout std_logic;
    bus11 : inout std_logic;
    bus12 : inout std_logic;
    bus13 : inout std_logic;
    bus14 : inout std_logic;
    bus15 : inout std_logic;
    bus16 : inout std_logic;
    bus17 : inout std_logic;
    bus18 : inout std_logic;
    bus19 : inout std_logic;
    bus2 : inout std_logic;
    bus20 : inout std_logic;
    bus21 : inout std_logic;
    bus22 : inout std_logic;
    bus23 : inout std_logic;
    bus24 : inout std_logic;
    bus25 : inout std_logic;
    bus26 : inout std_logic;
    bus27 : inout std_logic;
    bus28 : inout std_logic;
    bus29 : inout std_logic;
    bus3 : inout std_logic;
    bus30 : inout std_logic;
    bus31 : inout std_logic;
    bus4 : inout std_logic;
    bus5 : inout std_logic;
    bus6 : inout std_logic;
    bus7 : inout std_logic;
    bus8 : inout std_logic;
    bus9 : inout std_logic;
    \xbus ignpar in\ : inout std_logic;
    \xbus par in\ : inout std_logic;
    \xbus par out\ : inout std_logic;
    xdi0 : inout std_logic;
    xdi1 : inout std_logic;
    xdi10 : inout std_logic;
    xdi11 : inout std_logic;
    xdi12 : inout std_logic;
    xdi13 : inout std_logic;
    xdi14 : inout std_logic;
    xdi15 : inout std_logic;
    xdi16 : inout std_logic;
    xdi17 : inout std_logic;
    xdi18 : inout std_logic;
    xdi19 : inout std_logic;
    xdi2 : inout std_logic;
    xdi20 : inout std_logic;
    xdi21 : inout std_logic;
    xdi22 : inout std_logic;
    xdi23 : inout std_logic;
    xdi24 : inout std_logic;
    xdi25 : inout std_logic;
    xdi26 : inout std_logic;
    xdi27 : inout std_logic;
    xdi28 : inout std_logic;
    xdi29 : inout std_logic;
    xdi3 : inout std_logic;
    xdi30 : inout std_logic;
    xdi31 : inout std_logic;
    xdi4 : inout std_logic;
    xdi5 : inout std_logic;
    xdi6 : inout std_logic;
    xdi7 : inout std_logic;
    xdi8 : inout std_logic;
    xdi9 : inout std_logic;
    \hi 15-30\ : in std_logic
  );
end entity;
