library ieee;
use ieee.std_logic_1164.all;

package pages is

  component cadr4_clock1 is
    port (
      \-clock_reset_b\ : in std_logic;
      \-hang\ : in std_logic;
      \-ilong\ : in std_logic;
      \-tpdone\ : in std_logic;
      \-tpr0\ : out std_logic;
      \-tpr100\ : out std_logic;
      \-tpr105\ : out std_logic;
      \-tpr10\ : out std_logic;
      \-tpr110\ : out std_logic;
      \-tpr115\ : out std_logic;
      \-tpr120\ : out std_logic;
      \-tpr120a\ : out std_logic;
      \-tpr125\ : out std_logic;
      \-tpr140\ : out std_logic;
      \-tpr15\ : out std_logic;
      \-tpr160\ : out std_logic;
      \-tpr180\ : out std_logic;
      \-tpr200\ : out std_logic;
      \-tpr20\ : out std_logic;
      \-tpr20a\ : out std_logic;
      \-tpr25\ : out std_logic;
      \-tpr40\ : out std_logic;
      \-tpr5\ : out std_logic;
      \-tpr60\ : out std_logic;
      \-tpr65\ : out std_logic;
      \-tpr70\ : out std_logic;
      \-tpr75\ : out std_logic;
      \-tpr80\ : out std_logic;
      \-tpr80a\ : out std_logic;
      \-tpr85\ : out std_logic;
      \-tprend\ : out std_logic;
      \-tpw10\ : out std_logic;
      \-tpw20\ : out std_logic;
      \-tpw25\ : out std_logic;
      \-tpw30\ : out std_logic;
      \-tpw30a\ : out std_logic;
      \-tpw35\ : out std_logic;
      \-tpw40\ : out std_logic;
      \-tpw40a\ : out std_logic;
      \-tpw45\ : out std_logic;
      \-tpw50\ : out std_logic;
      \-tpw55\ : out std_logic;
      \-tpw60\ : out std_logic;
      \-tpw65\ : out std_logic;
      \-tpw70\ : out std_logic;
      \-tpw75\ : out std_logic;
      cyclecompleted : out std_logic;
      gnd : in std_logic;
      sspeed0 : in std_logic;
      sspeed1 : in std_logic;
      tprend : out std_logic
      );
  end component;

component cadr4_clock1 is
  port (
    \-destimod0\  : in std_logic;
    \-destimod1\  : in std_logic;
    \-destintctl\ : in std_logic;
    \-destlc\     : in std_logic;
    \-destmdr\    : in std_logic;
    \-destmem\    : in std_logic;
    \-destpdl(p)\ : in std_logic;
    \-destpdl(x)\ : in std_logic;
    \-destpdlp\   : in std_logic;
    \-destpdltop\ : in std_logic;
    \-destpdlx\   : in std_logic;
    \-destspc\    : in std_logic;
    \-destvma\    : in std_logic;
    \-div\        : in std_logic;
    \-funct0\     : in std_logic;
    \-funct1\     : in std_logic;
    \-funct2\     : in std_logic;
    \-funct3\     : in std_logic;
    \-idebug\     : in std_logic;
    \-ir22\       : in std_logic;
    \-ir25\       : in std_logic;
    \-ir31\       : in std_logic;
    \-iralu\      : in std_logic;
    \-irbyte\     : in std_logic;
    \-irdisp\     : in std_logic;
    \-irjump\     : in std_logic;
    \-mul\        : in std_logic;
    \-specalu\    : in std_logic;
    \-srcdc\      : in std_logic;
    \-srclc\      : in std_logic;
    \-srcmap\     : in std_logic;
    \-srcmd\      : in std_logic;
    \-srcopc\     : in std_logic;
    \-srcpdlidx\  : in std_logic;
    \-srcpdlpop\  : in std_logic;
    \-srcpdlptr\  : in std_logic;
    \-srcpdltop\  : in std_logic;
    \-srcq\       : in std_logic;
    \-srcspc\     : in std_logic;
    \-srcspcpop\  : in std_logic;
    \-srcvma\     : in std_logic;
    \destimod0_l\ : in std_logic;
    \iwrited_l\   : in std_logic;
    dest          : in std_logic;
    destm         : in std_logic;
    gnd           : in std_logic;
    hi5           : in std_logic;
    imod          : in std_logic;
    ir            : in std_logic_vector(0 to 48);
    iralu         : in std_logic;
    irdisp        : in std_logic;
    irjump        : in std_logic;
    nc            : in std_logic_vector(0 to 500)  -- Not connected ...
    );
end component;

end package;
