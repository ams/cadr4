library ieee;
use ieee.std_logic_1164.all;

entity cadr_mo1 is
  port (
    alu31  : in  std_logic;
    r31    : in  std_logic;
    a31b   : in  std_logic;
    ob31   : out std_logic;
    gnd    : in  std_logic;
    osel1a : in  std_logic;
    osel0a : in  std_logic;
    msk31  : in  std_logic;
    alu30  : in  std_logic;
    alu32  : in  std_logic;
    r30    : in  std_logic;
    a30    : in  std_logic;
    ob30   : out std_logic;
    msk30  : in  std_logic;
    alu29  : in  std_logic;
    r29    : in  std_logic;
    a29    : in  std_logic;
    ob29   : out std_logic;
    msk29  : in  std_logic;
    alu28  : in  std_logic;
    r28    : in  std_logic;
    a28    : in  std_logic;
    ob28   : out std_logic;
    msk28  : in  std_logic;
    alu27  : in  std_logic;
    alu23  : in  std_logic;
    r23    : in  std_logic;
    a23    : in  std_logic;
    ob23   : out std_logic;
    msk23  : in  std_logic;
    alu22  : in  std_logic;
    alu24  : in  std_logic;
    r22    : in  std_logic;
    a22    : in  std_logic;
    ob22   : out std_logic;
    msk22  : in  std_logic;
    alu21  : in  std_logic;
    r21    : in  std_logic;
    a21    : in  std_logic;
    ob21   : out std_logic;
    msk21  : in  std_logic;
    alu20  : in  std_logic;
    r20    : in  std_logic;
    a20    : in  std_logic;
    ob20   : out std_logic;
    msk20  : in  std_logic;
    alu19  : in  std_logic;
    r27    : in  std_logic;
    a27    : in  std_logic;
    ob27   : out std_logic;
    msk27  : in  std_logic;
    alu26  : in  std_logic;
    r24    : in  std_logic;
    a24    : in  std_logic;
    ob24   : out std_logic;
    msk24  : in  std_logic;
    alu25  : in  std_logic;
    r26    : in  std_logic;
    a26    : in  std_logic;
    ob26   : out std_logic;
    msk26  : in  std_logic;
    r25    : in  std_logic;
    a25    : in  std_logic;
    ob25   : out std_logic;
    msk25  : in  std_logic;
    r19    : in  std_logic;
    a19    : in  std_logic;
    ob19   : out std_logic;
    msk19  : in  std_logic;
    alu18  : in  std_logic;
    r18    : in  std_logic;
    a18    : in  std_logic;
    ob18   : out std_logic;
    msk18  : in  std_logic;
    r17    : in  std_logic;
    a17    : in  std_logic;
    ob17   : out std_logic;
    msk17  : in  std_logic;
    alu16  : in  std_logic;
    r16    : in  std_logic;
    a16    : in  std_logic;
    ob16   : out std_logic;
    msk16  : in  std_logic;
    alu15  : in  std_logic;
    alu17  : in  std_logic
    );
end;
