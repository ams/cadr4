-- The MIT CADR

library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;
use ttl.unsorted.all;

use work.utilities.all;

entity cadr4 is
end;

architecture structural of cadr4 is

  signal \-a31\                       : std_logic;
  signal \-aadr0a\                    : std_logic;
  signal \-aadr0b\                    : std_logic;
  signal \-aadr1a\                    : std_logic;
  signal \-aadr1b\                    : std_logic;
  signal \-aadr2a\                    : std_logic;
  signal \-aadr2b\                    : std_logic;
  signal \-aadr3a\                    : std_logic;
  signal \-aadr3b\                    : std_logic;
  signal \-aadr4a\                    : std_logic;
  signal \-aadr4b\                    : std_logic;
  signal \-aadr5a\                    : std_logic;
  signal \-aadr5b\                    : std_logic;
  signal \-aadr6a\                    : std_logic;
  signal \-aadr6b\                    : std_logic;
  signal \-aadr7a\                    : std_logic;
  signal \-aadr7b\                    : std_logic;
  signal \-aadr8a\                    : std_logic;
  signal \-aadr8b\                    : std_logic;
  signal \-aadr9a\                    : std_logic;
  signal \-aadr9b\                    : std_logic;
  signal \-adrpar\                    : std_logic;
  signal \-alu31\                     : std_logic;
  signal \-alu32\                     : std_logic;
  signal \-aluf0\                     : std_logic;
  signal \-aluf1\                     : std_logic;
  signal \-aluf2\                     : std_logic;
  signal \-aluf3\                     : std_logic;
  signal \-alumode\                   : std_logic;
  signal \-amemenb\                   : std_logic;
  signal \-apass\                     : std_logic;
  signal \-apassenb\                  : std_logic;
  signal \-ape\                       : std_logic;
  signal \-awpa\                      : std_logic;
  signal \-awpb\                      : std_logic;
  signal \-awpc\                      : std_logic;
  signal \-boot1\                     : std_logic;
  signal \-boot2\                     : std_logic;
  signal \-boot\                      : std_logic;
  signal \-bus.reset\                 : std_logic;
  signal \-busint.lm.reset\           : std_logic;
  signal \-cin0\                      : std_logic;
  signal \-cin12\                     : std_logic;
  signal \-cin16\                     : std_logic;
  signal \-cin20\                     : std_logic;
  signal \-cin24\                     : std_logic;
  signal \-cin28\                     : std_logic;
  signal \-cin32\                     : std_logic;
  signal \-cin4\                      : std_logic;
  signal \-cin8\                      : std_logic;
  signal \-clk0\                      : std_logic;
  signal \-clk1\                      : std_logic;
  signal \-clk2a\                     : std_logic;
  signal \-clk2c\                     : std_logic;
  signal \-clk3a\                     : std_logic;
  signal \-clk3d\                     : std_logic;
  signal \-clk3g\                     : std_logic;
  signal \-clk4a\                     : std_logic;
  signal \-clk4d\                     : std_logic;
  signal \-clk4e\                     : std_logic;
  signal \-clk5\                      : std_logic;
  signal \-clock_reset_a\             : std_logic;
  signal \-clock_reset_b\             : std_logic;
  signal \-dadr0a\                    : std_logic;
  signal \-dadr0b\                    : std_logic;
  signal \-dadr0c\                    : std_logic;
  signal \-dadr10a\                   : std_logic;
  signal \-dadr10c\                   : std_logic;
  signal \-dadr1a\                    : std_logic;
  signal \-dadr1b\                    : std_logic;
  signal \-dadr1c\                    : std_logic;
  signal \-dadr2a\                    : std_logic;
  signal \-dadr2b\                    : std_logic;
  signal \-dadr2c\                    : std_logic;
  signal \-dadr3a\                    : std_logic;
  signal \-dadr3b\                    : std_logic;
  signal \-dadr3c\                    : std_logic;
  signal \-dadr4a\                    : std_logic;
  signal \-dadr4b\                    : std_logic;
  signal \-dadr4c\                    : std_logic;
  signal \-dadr5a\                    : std_logic;
  signal \-dadr5b\                    : std_logic;
  signal \-dadr5c\                    : std_logic;
  signal \-dadr6a\                    : std_logic;
  signal \-dadr6b\                    : std_logic;
  signal \-dadr6c\                    : std_logic;
  signal \-dadr7a\                    : std_logic;
  signal \-dadr7b\                    : std_logic;
  signal \-dadr7c\                    : std_logic;
  signal \-dadr8a\                    : std_logic;
  signal \-dadr8b\                    : std_logic;
  signal \-dadr8c\                    : std_logic;
  signal \-dadr9a\                    : std_logic;
  signal \-dadr9b\                    : std_logic;
  signal \-dadr9c\                    : std_logic;
  signal \-dbread\                    : std_logic;
  signal \-dbwrite\                   : std_logic;
  signal \-destimod0\                 : std_logic;
  signal \-destimod1\                 : std_logic;
  signal \-destintctl\                : std_logic;
  signal \-destlc\                    : std_logic;
  signal \-destmdr\                   : std_logic;
  signal \-destmem\                   : std_logic;
  signal \-destpdl(p)\                : std_logic;
  signal \-destpdl(x)\                : std_logic;
  signal \-destpdlp\                  : std_logic;
  signal \-destpdltop\                : std_logic;
  signal \-destpdlx\                  : std_logic;
  signal \-destspc\                   : std_logic;
  signal \-destspcd\                  : std_logic;
  signal \-destvma\                   : std_logic;
  signal \-dfall\                     : std_logic;
  signal \-div\                       : std_logic;
  signal \-divposlasttime\            : std_logic;
  signal \-dmapbenb\                  : std_logic;
  signal \-dp\                        : std_logic;
  signal \-dparh\                     : std_logic;
  signal \-dpe\                       : std_logic;
  signal \-dr\                        : std_logic;
  signal \-dwea\                      : std_logic;
  signal \-dweb\                      : std_logic;
  signal \-dwec\                      : std_logic;
  signal \-errhalt\                   : std_logic;
  signal \-funct0\                    : std_logic;
  signal \-funct1\                    : std_logic;
  signal \-funct2\                    : std_logic;
  signal \-funct3\                    : std_logic;
  signal \-halt\                      : std_logic;
  signal \-halted\                    : std_logic;
  signal \-hang\                      : std_logic;
  signal \-higherr\                   : std_logic;
  signal \-ice0a\                     : std_logic;
  signal \-ice0b\                     : std_logic;
  signal \-ice0c\                     : std_logic;
  signal \-ice0d\                     : std_logic;
  signal \-ice1a\                     : std_logic;
  signal \-ice1b\                     : std_logic;
  signal \-ice1c\                     : std_logic;
  signal \-ice1d\                     : std_logic;
  signal \-ice2a\                     : std_logic;
  signal \-ice2b\                     : std_logic;
  signal \-ice2c\                     : std_logic;
  signal \-ice2d\                     : std_logic;
  signal \-ice3a\                     : std_logic;
  signal \-ice3b\                     : std_logic;
  signal \-ice3c\                     : std_logic;
  signal \-ice3d\                     : std_logic;
  signal \-idebug\                    : std_logic;
  signal \-ifetch\                    : std_logic;
  signal \-ignpar\                    : std_logic;
  signal \-ignpopj\                   : std_logic;
  signal \-ilong\                     : std_logic;
  signal \-imodd\                     : std_logic;
  signal \-inop\                      : std_logic;
  signal \-ipe\                       : std_logic;
  signal \-ipopj\                     : std_logic;
  signal \-ir0\                       : std_logic;
  signal \-ir12\                      : std_logic;
  signal \-ir13\                      : std_logic;
  signal \-ir1\                       : std_logic;
  signal \-ir22\                      : std_logic;
  signal \-ir25\                      : std_logic;
  signal \-ir2\                       : std_logic;
  signal \-ir31\                      : std_logic;
  signal \-ir3\                       : std_logic;
  signal \-ir4\                       : std_logic;
  signal \-ir6\                       : std_logic;
  signal \-ir8\                       : std_logic;
  signal \-iralu\                     : std_logic;
  signal \-irbyte\                    : std_logic;
  signal \-irdisp\                    : std_logic;
  signal \-irjump\                    : std_logic;
  signal \-iwea\                      : std_logic;
  signal \-iweb\                      : std_logic;
  signal \-iwec\                      : std_logic;
  signal \-iwed\                      : std_logic;
  signal \-iwee\                      : std_logic;
  signal \-iwef\                      : std_logic;
  signal \-iweg\                      : std_logic;
  signal \-iweh\                      : std_logic;
  signal \-iwei\                      : std_logic;
  signal \-iwej\                      : std_logic;
  signal \-iwek\                      : std_logic;
  signal \-iwel\                      : std_logic;
  signal \-iwem\                      : std_logic;
  signal \-iwen\                      : std_logic;
  signal \-iweo\                      : std_logic;
  signal \-iwep\                      : std_logic;
  signal \-iwrited\                   : std_logic;
  signal \-iwriteda\                  : std_logic;
  signal \-jcond\                     : std_logic;
  signal \-lc_modifies_mrot\          : std_logic;
  signal \-lcdrive\                   : std_logic;
  signal \-lcinc\                     : std_logic;
  signal \-lcry11\                    : std_logic;
  signal \-lcry15\                    : std_logic;
  signal \-lcry19\                    : std_logic;
  signal \-lcry23\                    : std_logic;
  signal \-lcry3\                     : std_logic;
  signal \-lcry7\                     : std_logic;
  signal \-ldclk\                     : std_logic;
  signal \-lddbirh\                   : std_logic;
  signal \-lddbirl\                   : std_logic;
  signal \-lddbirm\                   : std_logic;
  signal \-ldmode\                    : std_logic;
  signal \-ldopc\                     : std_logic;
  signal \-ldstat\                    : std_logic;
  signal \-loadmd\                    : std_logic;
  signal \-lowerhighok\               : std_logic;
  signal \-lparity\                   : std_logic;
  signal \-lparm\                     : std_logic;
  signal \-lpc.hold\                  : std_logic;
  signal \-lvmo22\                    : std_logic;
  signal \-lvmo23\                    : std_logic;
  signal \-machrun\                   : std_logic;
  signal \-machruna\                  : std_logic;
  signal \-madr0a\                    : std_logic;
  signal \-madr0b\                    : std_logic;
  signal \-madr1a\                    : std_logic;
  signal \-madr1b\                    : std_logic;
  signal \-madr2a\                    : std_logic;
  signal \-madr2b\                    : std_logic;
  signal \-madr3a\                    : std_logic;
  signal \-madr3b\                    : std_logic;
  signal \-madr4a\                    : std_logic;
  signal \-madr4b\                    : std_logic;
  signal \-mapdrive\                  : std_logic;
  signal \-mapi10a\                   : std_logic;
  signal \-mapi10b\                   : std_logic;
  signal \-mapi11a\                   : std_logic;
  signal \-mapi11b\                   : std_logic;
  signal \-mapi12a\                   : std_logic;
  signal \-mapi12b\                   : std_logic;
  signal \-mapi23\                    : std_logic;
  signal \-mapi8a\                    : std_logic;
  signal \-mapi8b\                    : std_logic;
  signal \-mapi9a\                    : std_logic;
  signal \-mapi9b\                    : std_logic;
  signal \-mbusy.sync\                : std_logic;
  signal \-mclk0\                     : std_logic;
  signal \-mclk1\                     : std_logic;
  signal \-mclk5\                     : std_logic;
  signal \-md0\                       : std_logic;
  signal \-md10\                      : std_logic;
  signal \-md11\                      : std_logic;
  signal \-md12\                      : std_logic;
  signal \-md13\                      : std_logic;
  signal \-md14\                      : std_logic;
  signal \-md15\                      : std_logic;
  signal \-md16\                      : std_logic;
  signal \-md17\                      : std_logic;
  signal \-md18\                      : std_logic;
  signal \-md19\                      : std_logic;
  signal \-md1\                       : std_logic;
  signal \-md20\                      : std_logic;
  signal \-md21\                      : std_logic;
  signal \-md22\                      : std_logic;
  signal \-md23\                      : std_logic;
  signal \-md24\                      : std_logic;
  signal \-md25\                      : std_logic;
  signal \-md26\                      : std_logic;
  signal \-md27\                      : std_logic;
  signal \-md28\                      : std_logic;
  signal \-md29\                      : std_logic;
  signal \-md2\                       : std_logic;
  signal \-md30\                      : std_logic;
  signal \-md31\                      : std_logic;
  signal \-md3\                       : std_logic;
  signal \-md4\                       : std_logic;
  signal \-md5\                       : std_logic;
  signal \-md6\                       : std_logic;
  signal \-md7\                       : std_logic;
  signal \-md8\                       : std_logic;
  signal \-md9\                       : std_logic;
  signal \-mddrive\                   : std_logic;
  signal \-mds0\                      : std_logic;
  signal \-mds10\                     : std_logic;
  signal \-mds11\                     : std_logic;
  signal \-mds12\                     : std_logic;
  signal \-mds13\                     : std_logic;
  signal \-mds14\                     : std_logic;
  signal \-mds15\                     : std_logic;
  signal \-mds16\                     : std_logic;
  signal \-mds17\                     : std_logic;
  signal \-mds18\                     : std_logic;
  signal \-mds19\                     : std_logic;
  signal \-mds1\                      : std_logic;
  signal \-mds20\                     : std_logic;
  signal \-mds21\                     : std_logic;
  signal \-mds22\                     : std_logic;
  signal \-mds23\                     : std_logic;
  signal \-mds24\                     : std_logic;
  signal \-mds25\                     : std_logic;
  signal \-mds26\                     : std_logic;
  signal \-mds27\                     : std_logic;
  signal \-mds28\                     : std_logic;
  signal \-mds29\                     : std_logic;
  signal \-mds2\                      : std_logic;
  signal \-mds30\                     : std_logic;
  signal \-mds31\                     : std_logic;
  signal \-mds3\                      : std_logic;
  signal \-mds4\                      : std_logic;
  signal \-mds5\                      : std_logic;
  signal \-mds6\                      : std_logic;
  signal \-mds7\                      : std_logic;
  signal \-mds8\                      : std_logic;
  signal \-mds9\                      : std_logic;
  signal \-memack\                    : std_logic;
  signal \-memdrive.a\                : std_logic;
  signal \-memdrive.b\                : std_logic;
  signal \-memgrant\                  : std_logic;
  signal \-memop\                     : std_logic;
  signal \-memparok\                  : std_logic;
  signal \-mempe\                     : std_logic;
  signal \-memprepare\                : std_logic;
  signal \-memrd\                     : std_logic;
  signal \-memrq\                     : std_logic;
  signal \-memstart\                  : std_logic;
  signal \-memwr\                     : std_logic;
  signal \-mfdrive\                   : std_logic;
  signal \-mfinish\                   : std_logic;
  signal \-mfinishd\                  : std_logic;
  signal \-mpass\                     : std_logic;
  signal \-mpassl\                    : std_logic;
  signal \-mpassm\                    : std_logic;
  signal \-mpe\                       : std_logic;
  signal \-mr\                        : std_logic;
  signal \-mul\                       : std_logic;
  signal \-mulnop\                    : std_logic;
  signal \-mwpa\                      : std_logic;
  signal \-mwpb\                      : std_logic;
  signal \-needfetch\                 : std_logic;
  signal \-newlc.in\                  : std_logic;
  signal \-newlc\                     : std_logic;
  signal \-nop11\                     : std_logic;
  signal \-nop\                       : std_logic;
  signal \-nopa\                      : std_logic;
  signal \-opcclk\                    : std_logic;
  signal \-opcdrive\                  : std_logic;
  signal \-opcinh\                    : std_logic;
  signal \-parerr\                    : std_logic;
  signal \-pc12b\                     : std_logic;
  signal \-pc13b\                     : std_logic;
  signal \-pcb0\                      : std_logic;
  signal \-pcb10\                     : std_logic;
  signal \-pcb11\                     : std_logic;
  signal \-pcb1\                      : std_logic;
  signal \-pcb2\                      : std_logic;
  signal \-pcb3\                      : std_logic;
  signal \-pcb4\                      : std_logic;
  signal \-pcb5\                      : std_logic;
  signal \-pcb6\                      : std_logic;
  signal \-pcb7\                      : std_logic;
  signal \-pcb8\                      : std_logic;
  signal \-pcb9\                      : std_logic;
  signal \-pcc0\                      : std_logic;
  signal \-pcc10\                     : std_logic;
  signal \-pcc11\                     : std_logic;
  signal \-pcc1\                      : std_logic;
  signal \-pcc2\                      : std_logic;
  signal \-pcc3\                      : std_logic;
  signal \-pcc4\                      : std_logic;
  signal \-pcc5\                      : std_logic;
  signal \-pcc6\                      : std_logic;
  signal \-pcc7\                      : std_logic;
  signal \-pcc8\                      : std_logic;
  signal \-pcc9\                      : std_logic;
  signal \-pdla0a\                    : std_logic;
  signal \-pdla0b\                    : std_logic;
  signal \-pdla1a\                    : std_logic;
  signal \-pdla1b\                    : std_logic;
  signal \-pdla2a\                    : std_logic;
  signal \-pdla2b\                    : std_logic;
  signal \-pdla3a\                    : std_logic;
  signal \-pdla3b\                    : std_logic;
  signal \-pdla4a\                    : std_logic;
  signal \-pdla4b\                    : std_logic;
  signal \-pdla5a\                    : std_logic;
  signal \-pdla5b\                    : std_logic;
  signal \-pdla6a\                    : std_logic;
  signal \-pdla6b\                    : std_logic;
  signal \-pdla7a\                    : std_logic;
  signal \-pdla7b\                    : std_logic;
  signal \-pdla8a\                    : std_logic;
  signal \-pdla8b\                    : std_logic;
  signal \-pdla9a\                    : std_logic;
  signal \-pdla9b\                    : std_logic;
  signal \-pdlcnt\                    : std_logic;
  signal \-pdlcry3\                   : std_logic;
  signal \-pdlcry7\                   : std_logic;
  signal \-pdldrive\                  : std_logic;
  signal \-pdlpa\                     : std_logic;
  signal \-pdlpb\                     : std_logic;
  signal \-pdlpe\                     : std_logic;
  signal \-pdlwrited\                 : std_logic;
  signal \-pfr\                       : std_logic;
  signal \-pfw\                       : std_logic;
  signal \-pma10\                     : std_logic;
  signal \-pma11\                     : std_logic;
  signal \-pma12\                     : std_logic;
  signal \-pma13\                     : std_logic;
  signal \-pma14\                     : std_logic;
  signal \-pma15\                     : std_logic;
  signal \-pma16\                     : std_logic;
  signal \-pma17\                     : std_logic;
  signal \-pma18\                     : std_logic;
  signal \-pma19\                     : std_logic;
  signal \-pma20\                     : std_logic;
  signal \-pma21\                     : std_logic;
  signal \-pma8\                      : std_logic;
  signal \-pma9\                      : std_logic;
  signal \-popj\                      : std_logic;
  signal \-power_reset\               : std_logic;
  signal \-ppdrive\                   : std_logic;
  signal \-prog.reset\                : std_logic;
  signal \-promce0\                   : std_logic;
  signal \-promce1\                   : std_logic;
  signal \-promdisabled\              : std_logic;
  signal \-promenable\                : std_logic;
  signal \-prompc0\                   : std_logic;
  signal \-prompc1\                   : std_logic;
  signal \-prompc2\                   : std_logic;
  signal \-prompc3\                   : std_logic;
  signal \-prompc4\                   : std_logic;
  signal \-prompc5\                   : std_logic;
  signal \-prompc6\                   : std_logic;
  signal \-prompc7\                   : std_logic;
  signal \-prompc8\                   : std_logic;
  signal \-prompc9\                   : std_logic;
  signal \-pwidx\                     : std_logic;
  signal \-pwpa\                      : std_logic;
  signal \-pwpb\                      : std_logic;
  signal \-pwpc\                      : std_logic;
  signal \-qdrive\                    : std_logic;
  signal \-rdfinish\                  : std_logic;
  signal \-reset\                     : std_logic;
  signal \-run\                       : std_logic;
  signal \-s4\                        : std_logic;
  signal \-sh3\                       : std_logic;
  signal \-sh4\                       : std_logic;
  signal \-spccry\                    : std_logic;
  signal \-spcdrive\                  : std_logic;
  signal \-spcnt\                     : std_logic;
  signal \-spcpass\                   : std_logic;
  signal \-spcwparl\                  : std_logic;
  signal \-spcwpass\                  : std_logic;
  signal \-spe\                       : std_logic;
  signal \-specalu\                   : std_logic;
  signal \-spop\                      : std_logic;
  signal \-spush\                     : std_logic;
  signal \-spushd\                    : std_logic;
  signal \-spy.ah\                    : std_logic;
  signal \-spy.al\                    : std_logic;
  signal \-spy.flag1\                 : std_logic;
  signal \-spy.flag2\                 : std_logic;
  signal \-spy.irh\                   : std_logic;
  signal \-spy.irl\                   : std_logic;
  signal \-spy.irm\                   : std_logic;
  signal \-spy.mh\                    : std_logic;
  signal \-spy.ml\                    : std_logic;
  signal \-spy.obh\                   : std_logic;
  signal \-spy.obl\                   : std_logic;
  signal \-spy.opc\                   : std_logic;
  signal \-spy.pc\                    : std_logic;
  signal \-spy.sth\                   : std_logic;
  signal \-spy.stl\                   : std_logic;
  signal \-sr\                        : std_logic;
  signal \-srcdc\                     : std_logic;
  signal \-srclc\                     : std_logic;
  signal \-srcm\                      : std_logic;
  signal \-srcmap\                    : std_logic;
  signal \-srcmd\                     : std_logic;
  signal \-srcopc\                    : std_logic;
  signal \-srcpdlidx\                 : std_logic;
  signal \-srcpdlpop\                 : std_logic;
  signal \-srcpdlptr\                 : std_logic;
  signal \-srcpdltop\                 : std_logic;
  signal \-srcq\                      : std_logic;
  signal \-srcspc\                    : std_logic;
  signal \-srcspcpop\                 : std_logic;
  signal \-srcspcpopreal\             : std_logic;
  signal \-srcvma\                    : std_logic;
  signal \-ssdone\                    : std_logic;
  signal \-statbit\                   : std_logic;
  signal \-stathalt\                  : std_logic;
  signal \-stc12\                     : std_logic;
  signal \-stc16\                     : std_logic;
  signal \-stc20\                     : std_logic;
  signal \-stc24\                     : std_logic;
  signal \-stc28\                     : std_logic;
  signal \-stc32\                     : std_logic;
  signal \-stc4\                      : std_logic;
  signal \-stc8\                      : std_logic;
  signal \-step\                      : std_logic;
  signal \-swpa\                      : std_logic;
  signal \-swpb\                      : std_logic;
  signal \-tpclk\                     : std_logic;
  signal \-tpdone\                    : std_logic;
  signal \-tpr0\                      : std_logic;
  signal \-tpr100\                    : std_logic;
  signal \-tpr105\                    : std_logic;
  signal \-tpr10\                     : std_logic;
  signal \-tpr110\                    : std_logic;
  signal \-tpr115\                    : std_logic;
  signal \-tpr120\                    : std_logic;
  signal \-tpr120a\                   : std_logic;
  signal \-tpr125\                    : std_logic;
  signal \-tpr140\                    : std_logic;
  signal \-tpr15\                     : std_logic;
  signal \-tpr160\                    : std_logic;
  signal \-tpr180\                    : std_logic;
  signal \-tpr200\                    : std_logic;
  signal \-tpr20\                     : std_logic;
  signal \-tpr20a\                    : std_logic;
  signal \-tpr25\                     : std_logic;
  signal \-tpr40\                     : std_logic;
  signal \-tpr5\                      : std_logic;
  signal \-tpr60\                     : std_logic;
  signal \-tpr65\                     : std_logic;
  signal \-tpr70\                     : std_logic;
  signal \-tpr75\                     : std_logic;
  signal \-tpr80\                     : std_logic;
  signal \-tpr80a\                    : std_logic;
  signal \-tpr85\                     : std_logic;
  signal \-tprend\                    : std_logic;
  signal \-tptse\                     : std_logic;
  signal \-tpw10\                     : std_logic;
  signal \-tpw20\                     : std_logic;
  signal \-tpw25\                     : std_logic;
  signal \-tpw30\                     : std_logic;
  signal \-tpw30a\                    : std_logic;
  signal \-tpw35\                     : std_logic;
  signal \-tpw40\                     : std_logic;
  signal \-tpw40a\                    : std_logic;
  signal \-tpw45\                     : std_logic;
  signal \-tpw50\                     : std_logic;
  signal \-tpw55\                     : std_logic;
  signal \-tpw60\                     : std_logic;
  signal \-tpw65\                     : std_logic;
  signal \-tpw70\                     : std_logic;
  signal \-tpw75\                     : std_logic;
  signal \-trap\                      : std_logic;
  signal \-trapenb\                   : std_logic;
  signal \-tse1\                      : std_logic;
  signal \-tse2\                      : std_logic;
  signal \-tse3\                      : std_logic;
  signal \-tse4\                      : std_logic;
  signal \-upperhighok\               : std_logic;
  signal \-use.map\                   : std_logic;
  signal \-v0pe\                      : std_logic;
  signal \-v1pe\                      : std_logic;
  signal \-vm0wpa\                    : std_logic;
  signal \-vm0wpb\                    : std_logic;
  signal \-vm1lpar\                   : std_logic;
  signal \-vm1wpa\                    : std_logic;
  signal \-vm1wpb\                    : std_logic;
  signal \-vma0\                      : std_logic;
  signal \-vma10\                     : std_logic;
  signal \-vma11\                     : std_logic;
  signal \-vma12\                     : std_logic;
  signal \-vma13\                     : std_logic;
  signal \-vma14\                     : std_logic;
  signal \-vma15\                     : std_logic;
  signal \-vma16\                     : std_logic;
  signal \-vma17\                     : std_logic;
  signal \-vma18\                     : std_logic;
  signal \-vma19\                     : std_logic;
  signal \-vma1\                      : std_logic;
  signal \-vma20\                     : std_logic;
  signal \-vma21\                     : std_logic;
  signal \-vma22\                     : std_logic;
  signal \-vma23\                     : std_logic;
  signal \-vma24\                     : std_logic;
  signal \-vma25\                     : std_logic;
  signal \-vma26\                     : std_logic;
  signal \-vma27\                     : std_logic;
  signal \-vma28\                     : std_logic;
  signal \-vma29\                     : std_logic;
  signal \-vma2\                      : std_logic;
  signal \-vma30\                     : std_logic;
  signal \-vma31\                     : std_logic;
  signal \-vma3\                      : std_logic;
  signal \-vma4\                      : std_logic;
  signal \-vma5\                      : std_logic;
  signal \-vma6\                      : std_logic;
  signal \-vma7\                      : std_logic;
  signal \-vma8\                      : std_logic;
  signal \-vma9\                      : std_logic;
  signal \-vmadrive\                  : std_logic;
  signal \-vmaenb\                    : std_logic;
  signal \-vmaok\                     : std_logic;
  signal \-vmap0\                     : std_logic;
  signal \-vmap1\                     : std_logic;
  signal \-vmap2\                     : std_logic;
  signal \-vmap3\                     : std_logic;
  signal \-vmap4\                     : std_logic;
  signal \-vmas0\                     : std_logic;
  signal \-vmas10\                    : std_logic;
  signal \-vmas11\                    : std_logic;
  signal \-vmas12\                    : std_logic;
  signal \-vmas13\                    : std_logic;
  signal \-vmas14\                    : std_logic;
  signal \-vmas15\                    : std_logic;
  signal \-vmas16\                    : std_logic;
  signal \-vmas17\                    : std_logic;
  signal \-vmas18\                    : std_logic;
  signal \-vmas19\                    : std_logic;
  signal \-vmas1\                     : std_logic;
  signal \-vmas20\                    : std_logic;
  signal \-vmas21\                    : std_logic;
  signal \-vmas22\                    : std_logic;
  signal \-vmas23\                    : std_logic;
  signal \-vmas24\                    : std_logic;
  signal \-vmas25\                    : std_logic;
  signal \-vmas26\                    : std_logic;
  signal \-vmas27\                    : std_logic;
  signal \-vmas28\                    : std_logic;
  signal \-vmas29\                    : std_logic;
  signal \-vmas2\                     : std_logic;
  signal \-vmas30\                    : std_logic;
  signal \-vmas31\                    : std_logic;
  signal \-vmas3\                     : std_logic;
  signal \-vmas4\                     : std_logic;
  signal \-vmas5\                     : std_logic;
  signal \-vmas6\                     : std_logic;
  signal \-vmas7\                     : std_logic;
  signal \-vmas8\                     : std_logic;
  signal \-vmas9\                     : std_logic;
  signal \-vmo0\                      : std_logic;
  signal \-vmo10\                     : std_logic;
  signal \-vmo11\                     : std_logic;
  signal \-vmo12\                     : std_logic;
  signal \-vmo13\                     : std_logic;
  signal \-vmo14\                     : std_logic;
  signal \-vmo15\                     : std_logic;
  signal \-vmo16\                     : std_logic;
  signal \-vmo17\                     : std_logic;
  signal \-vmo18\                     : std_logic;
  signal \-vmo19\                     : std_logic;
  signal \-vmo1\                      : std_logic;
  signal \-vmo20\                     : std_logic;
  signal \-vmo21\                     : std_logic;
  signal \-vmo22\                     : std_logic;
  signal \-vmo23\                     : std_logic;
  signal \-vmo2\                      : std_logic;
  signal \-vmo3\                      : std_logic;
  signal \-vmo4\                      : std_logic;
  signal \-vmo5\                      : std_logic;
  signal \-vmo6\                      : std_logic;
  signal \-vmo7\                      : std_logic;
  signal \-vmo8\                      : std_logic;
  signal \-vmo9\                      : std_logic;
  signal \-wait\                      : std_logic;
  signal \-wmap\                      : std_logic;
  signal \-wmapd\                     : std_logic;
  signal \-wp1\                       : std_logic;
  signal \-wp2\                       : std_logic;
  signal \-wp3\                       : std_logic;
  signal \-wp4\                       : std_logic;
  signal \-wp5\                       : std_logic;
  signal \-zero16.drive\              : std_logic;
  signal \boot.trap\                  : std_logic;
  signal \bottom.1k\                  : std_logic;
  signal \bus.power.reset_l\          : std_logic;
  signal \destimod0_l\                : std_logic;
  signal \have_wrong_word\            : std_logic;
  signal \inst_in_2nd_or_4th_quarter\ : std_logic;
  signal \inst_in_left_half\          : std_logic;
  signal \int.enable\                 : std_logic;
  signal \iwrited_l\                  : std_logic;
  signal \last_byte_in_word\          : std_logic;
  signal \lc_byte_mode\               : std_logic;
  signal \lm_drive_enb\               : std_logic;
  signal \lpc.hold\                   : std_logic;
  signal \machruna_l\                 : std_logic;
  signal \mbusy.sync\                 : std_logic;
  signal \mempar_in\                  : std_logic;
  signal \mempar_out\                 : std_logic;
  signal \next.instr\                 : std_logic;
  signal \next.instrd\                : std_logic;
  signal \pgf.or.int.or.sb\           : std_logic;
  signal \pgf.or.int\                 : std_logic;
  signal \power_reset_a\              : std_logic;
  signal \prog.boot\                  : std_logic;
  signal \prog.bus.reset\             : std_logic;
  signal \prog.unibus.reset\          : std_logic;
  signal \rd.in.progress\             : std_logic;
  signal \sequence.break\             : std_logic;
  signal \set.rd.in.progress\         : std_logic;
  signal \stat.ovf\                   : std_logic;
  signal \use.md\                     : std_logic;
  signal \zero12.drive\               : std_logic;
  signal \zero16.drive\               : std_logic;
  signal a0                           : std_logic;
  signal a10                          : std_logic;
  signal a11                          : std_logic;
  signal a12                          : std_logic;
  signal a13                          : std_logic;
  signal a14                          : std_logic;
  signal a15                          : std_logic;
  signal a16                          : std_logic;
  signal a17                          : std_logic;
  signal a18                          : std_logic;
  signal a19                          : std_logic;
  signal a1                           : std_logic;
  signal a20                          : std_logic;
  signal a21                          : std_logic;
  signal a22                          : std_logic;
  signal a23                          : std_logic;
  signal a24                          : std_logic;
  signal a25                          : std_logic;
  signal a26                          : std_logic;
  signal a27                          : std_logic;
  signal a28                          : std_logic;
  signal a29                          : std_logic;
  signal a2                           : std_logic;
  signal a30                          : std_logic;
  signal a31a                         : std_logic;
  signal a31b                         : std_logic;
  signal a3                           : std_logic;
  signal a4                           : std_logic;
  signal a5                           : std_logic;
  signal a6                           : std_logic;
  signal a7                           : std_logic;
  signal a8                           : std_logic;
  signal a9                           : std_logic;
  signal aa0                          : std_logic;
  signal aa10                         : std_logic;
  signal aa11                         : std_logic;
  signal aa12                         : std_logic;
  signal aa13                         : std_logic;
  signal aa14                         : std_logic;
  signal aa15                         : std_logic;
  signal aa16                         : std_logic;
  signal aa17                         : std_logic;
  signal aa1                          : std_logic;
  signal aa2                          : std_logic;
  signal aa3                          : std_logic;
  signal aa4                          : std_logic;
  signal aa5                          : std_logic;
  signal aa6                          : std_logic;
  signal aa7                          : std_logic;
  signal aa8                          : std_logic;
  signal aa9                          : std_logic;
  signal aeqm                         : std_logic;
  signal alu0                         : std_logic;
  signal alu10                        : std_logic;
  signal alu11                        : std_logic;
  signal alu12                        : std_logic;
  signal alu13                        : std_logic;
  signal alu14                        : std_logic;
  signal alu15                        : std_logic;
  signal alu16                        : std_logic;
  signal alu17                        : std_logic;
  signal alu18                        : std_logic;
  signal alu19                        : std_logic;
  signal alu1                         : std_logic;
  signal alu20                        : std_logic;
  signal alu21                        : std_logic;
  signal alu22                        : std_logic;
  signal alu23                        : std_logic;
  signal alu24                        : std_logic;
  signal alu25                        : std_logic;
  signal alu26                        : std_logic;
  signal alu27                        : std_logic;
  signal alu28                        : std_logic;
  signal alu29                        : std_logic;
  signal alu2                         : std_logic;
  signal alu30                        : std_logic;
  signal alu31                        : std_logic;
  signal alu32                        : std_logic;
  signal alu3                         : std_logic;
  signal alu4                         : std_logic;
  signal alu5                         : std_logic;
  signal alu6                         : std_logic;
  signal alu7                         : std_logic;
  signal alu8                         : std_logic;
  signal alu9                         : std_logic;
  signal aluadd                       : std_logic;
  signal aluf0a                       : std_logic;
  signal aluf0b                       : std_logic;
  signal aluf1a                       : std_logic;
  signal aluf1b                       : std_logic;
  signal aluf2a                       : std_logic;
  signal aluf2b                       : std_logic;
  signal aluf3a                       : std_logic;
  signal aluf3b                       : std_logic;
  signal alumode                      : std_logic;
  signal aluneg                       : std_logic;
  signal alusub                       : std_logic;
  signal amem0                        : std_logic;
  signal amem10                       : std_logic;
  signal amem11                       : std_logic;
  signal amem12                       : std_logic;
  signal amem13                       : std_logic;
  signal amem14                       : std_logic;
  signal amem15                       : std_logic;
  signal amem16                       : std_logic;
  signal amem17                       : std_logic;
  signal amem18                       : std_logic;
  signal amem19                       : std_logic;
  signal amem1                        : std_logic;
  signal amem20                       : std_logic;
  signal amem21                       : std_logic;
  signal amem22                       : std_logic;
  signal amem23                       : std_logic;
  signal amem24                       : std_logic;
  signal amem25                       : std_logic;
  signal amem26                       : std_logic;
  signal amem27                       : std_logic;
  signal amem28                       : std_logic;
  signal amem29                       : std_logic;
  signal amem2                        : std_logic;
  signal amem30                       : std_logic;
  signal amem31                       : std_logic;
  signal amem3                        : std_logic;
  signal amem4                        : std_logic;
  signal amem5                        : std_logic;
  signal amem6                        : std_logic;
  signal amem7                        : std_logic;
  signal amem8                        : std_logic;
  signal amem9                        : std_logic;
  signal amemparity                   : std_logic;
  signal aparity                      : std_logic;
  signal aparl                        : std_logic;
  signal aparm                        : std_logic;
  signal aparok                       : std_logic;
  signal apass1                       : std_logic;
  signal apass2                       : std_logic;
  signal apassenb                     : std_logic;
  signal clk1                         : std_logic;
  signal clk1a                        : std_logic;
  signal clk2                         : std_logic;
  signal clk2a                        : std_logic;
  signal clk2b                        : std_logic;
  signal clk2c                        : std_logic;
  signal clk3                         : std_logic;
  signal clk3a                        : std_logic;
  signal clk3b                        : std_logic;
  signal clk3c                        : std_logic;
  signal clk3d                        : std_logic;
  signal clk3e                        : std_logic;
  signal clk3f                        : std_logic;
  signal clk4                         : std_logic;
  signal clk4a                        : std_logic;
  signal clk4b                        : std_logic;
  signal clk4c                        : std_logic;
  signal clk4d                        : std_logic;
  signal clk4e                        : std_logic;
  signal clk4f                        : std_logic;
  signal clk5                         : std_logic;
  signal clk5a                        : std_logic;
  signal conds0                       : std_logic;
  signal conds1                       : std_logic;
  signal conds2                       : std_logic;
  signal cyclecompleted               : std_logic;
  signal dadr10a                      : std_logic;
  signal dadr10c                      : std_logic;
  signal dc0                          : std_logic;
  signal dc1                          : std_logic;
  signal dc2                          : std_logic;
  signal dc3                          : std_logic;
  signal dc4                          : std_logic;
  signal dc5                          : std_logic;
  signal dc6                          : std_logic;
  signal dc7                          : std_logic;
  signal dc8                          : std_logic;
  signal dc9                          : std_logic;
  signal dcdrive                      : std_logic;
  signal dest                         : std_logic;
  signal destd                        : std_logic;
  signal destm                        : std_logic;
  signal destmd                       : std_logic;
  signal destmdr                      : std_logic;
  signal destmem                      : std_logic;
  signal destspc                      : std_logic;
  signal destspcd                     : std_logic;
  signal dispenb                      : std_logic;
  signal dispwr                       : std_logic;
  signal divaddcond                   : std_logic;
  signal divsubcond                   : std_logic;
  signal dmask0                       : std_logic;
  signal dmask1                       : std_logic;
  signal dmask2                       : std_logic;
  signal dmask3                       : std_logic;
  signal dmask4                       : std_logic;
  signal dmask5                       : std_logic;
  signal dmask6                       : std_logic;
  signal dn                           : std_logic;
  signal dp                           : std_logic;
  signal dpar                         : std_logic;
  signal dpareven                     : std_logic;
  signal dparl                        : std_logic;
  signal dparok                       : std_logic;
  signal dpc0                         : std_logic;
  signal dpc10                        : std_logic;
  signal dpc11                        : std_logic;
  signal dpc12                        : std_logic;
  signal dpc13                        : std_logic;
  signal dpc1                         : std_logic;
  signal dpc2                         : std_logic;
  signal dpc3                         : std_logic;
  signal dpc4                         : std_logic;
  signal dpc5                         : std_logic;
  signal dpc6                         : std_logic;
  signal dpc7                         : std_logic;
  signal dpc8                         : std_logic;
  signal dpc9                         : std_logic;
  signal dpe                          : std_logic;
  signal dr                           : std_logic;
  signal eadr0                        : std_logic;
  signal eadr1                        : std_logic;
  signal eadr2                        : std_logic;
  signal eadr3                        : std_logic;
  signal err                          : std_logic;
  signal errstop                      : std_logic;
  signal g2b                          : std_logic;
  signal gnd                          : std_logic;
  signal hi10                         : std_logic;
  signal hi11                         : std_logic;
  signal hi12                         : std_logic;
  signal hi1                          : std_logic;
  signal hi2                          : std_logic;
  signal hi3                          : std_logic;
  signal hi4                          : std_logic;
  signal hi5                          : std_logic;
  signal hi6                          : std_logic;
  signal hi7                          : std_logic;
  signal hi8                          : std_logic;
  signal hi9                          : std_logic;
  signal highok                       : std_logic;
  signal i0                           : std_logic;
  signal i10                          : std_logic;
  signal i11                          : std_logic;
  signal i12                          : std_logic;
  signal i13                          : std_logic;
  signal i14                          : std_logic;
  signal i15                          : std_logic;
  signal i16                          : std_logic;
  signal i17                          : std_logic;
  signal i18                          : std_logic;
  signal i19                          : std_logic;
  signal i1                           : std_logic;
  signal i20                          : std_logic;
  signal i21                          : std_logic;
  signal i22                          : std_logic;
  signal i23                          : std_logic;
  signal i24                          : std_logic;
  signal i25                          : std_logic;
  signal i26                          : std_logic;
  signal i27                          : std_logic;
  signal i28                          : std_logic;
  signal i29                          : std_logic;
  signal i2                           : std_logic;
  signal i30                          : std_logic;
  signal i31                          : std_logic;
  signal i32                          : std_logic;
  signal i33                          : std_logic;
  signal i34                          : std_logic;
  signal i35                          : std_logic;
  signal i36                          : std_logic;
  signal i37                          : std_logic;
  signal i38                          : std_logic;
  signal i39                          : std_logic;
  signal i3                           : std_logic;
  signal i40                          : std_logic;
  signal i41                          : std_logic;
  signal i42                          : std_logic;
  signal i43                          : std_logic;
  signal i44                          : std_logic;
  signal i45                          : std_logic;
  signal i46                          : std_logic;
  signal i47                          : std_logic;
  signal i48                          : std_logic;
  signal i4                           : std_logic;
  signal i5                           : std_logic;
  signal i6                           : std_logic;
  signal i7                           : std_logic;
  signal i8                           : std_logic;
  signal i9                           : std_logic;
  signal idebug                       : std_logic;
  signal imod                         : std_logic;
  signal imodd                        : std_logic;
  signal inop                         : std_logic;
  signal int                          : std_logic;
  signal internal10                   : std_logic;
  signal internal11                   : std_logic;
  signal internal12                   : std_logic;
  signal internal13                   : std_logic;
  signal internal14                   : std_logic;
  signal internal15                   : std_logic;
  signal internal16                   : std_logic;
  signal internal17                   : std_logic;
  signal internal18                   : std_logic;
  signal internal19                   : std_logic;
  signal internal1                    : std_logic;
  signal internal20                   : std_logic;
  signal internal21                   : std_logic;
  signal internal22                   : std_logic;
  signal internal23                   : std_logic;
  signal internal24                   : std_logic;
  signal internal25                   : std_logic;
  signal internal26                   : std_logic;
  signal internal27                   : std_logic;
  signal internal28                   : std_logic;
  signal internal29                   : std_logic;
  signal internal2                    : std_logic;
  signal internal30                   : std_logic;
  signal internal31                   : std_logic;
  signal internal32                   : std_logic;
  signal internal33                   : std_logic;
  signal internal34                   : std_logic;
  signal internal35                   : std_logic;
  signal internal36                   : std_logic;
  signal internal37                   : std_logic;
  signal internal3                    : std_logic;
  signal internal4                    : std_logic;
  signal internal5                    : std_logic;
  signal internal7                    : std_logic;
  signal internal8                    : std_logic;
  signal internal9                    : std_logic;
  signal iob0                         : std_logic;
  signal iob10                        : std_logic;
  signal iob11                        : std_logic;
  signal iob12                        : std_logic;
  signal iob13                        : std_logic;
  signal iob14                        : std_logic;
  signal iob15                        : std_logic;
  signal iob16                        : std_logic;
  signal iob17                        : std_logic;
  signal iob18                        : std_logic;
  signal iob19                        : std_logic;
  signal iob1                         : std_logic;
  signal iob20                        : std_logic;
  signal iob21                        : std_logic;
  signal iob22                        : std_logic;
  signal iob23                        : std_logic;
  signal iob24                        : std_logic;
  signal iob25                        : std_logic;
  signal iob26                        : std_logic;
  signal iob27                        : std_logic;
  signal iob28                        : std_logic;
  signal iob29                        : std_logic;
  signal iob2                         : std_logic;
  signal iob30                        : std_logic;
  signal iob31                        : std_logic;
  signal iob32                        : std_logic;
  signal iob33                        : std_logic;
  signal iob34                        : std_logic;
  signal iob35                        : std_logic;
  signal iob36                        : std_logic;
  signal iob37                        : std_logic;
  signal iob38                        : std_logic;
  signal iob39                        : std_logic;
  signal iob3                         : std_logic;
  signal iob40                        : std_logic;
  signal iob41                        : std_logic;
  signal iob42                        : std_logic;
  signal iob43                        : std_logic;
  signal iob44                        : std_logic;
  signal iob45                        : std_logic;
  signal iob46                        : std_logic;
  signal iob47                        : std_logic;
  signal iob4                         : std_logic;
  signal iob5                         : std_logic;
  signal iob6                         : std_logic;
  signal iob7                         : std_logic;
  signal iob8                         : std_logic;
  signal iob9                         : std_logic;
  signal ipar0                        : std_logic;
  signal ipar1                        : std_logic;
  signal ipar2                        : std_logic;
  signal ipar3                        : std_logic;
  signal iparity                      : std_logic;
  signal iparok                       : std_logic;
  signal ipc0                         : std_logic;
  signal ipc10                        : std_logic;
  signal ipc11                        : std_logic;
  signal ipc12                        : std_logic;
  signal ipc13                        : std_logic;
  signal ipc1                         : std_logic;
  signal ipc2                         : std_logic;
  signal ipc3                         : std_logic;
  signal ipc4                         : std_logic;
  signal ipc5                         : std_logic;
  signal ipc6                         : std_logic;
  signal ipc7                         : std_logic;
  signal ipc8                         : std_logic;
  signal ipc9                         : std_logic;
  signal ipe                          : std_logic;
  signal ir0                          : std_logic;
  signal ir10                         : std_logic;
  signal ir11                         : std_logic;
  signal ir12                         : std_logic;
  signal ir12b                        : std_logic;
  signal ir13                         : std_logic;
  signal ir13b                        : std_logic;
  signal ir14                         : std_logic;
  signal ir14b                        : std_logic;
  signal ir15                         : std_logic;
  signal ir15b                        : std_logic;
  signal ir16                         : std_logic;
  signal ir16b                        : std_logic;
  signal ir17                         : std_logic;
  signal ir17b                        : std_logic;
  signal ir18                         : std_logic;
  signal ir18b                        : std_logic;
  signal ir19                         : std_logic;
  signal ir19b                        : std_logic;
  signal ir1                          : std_logic;
  signal ir20                         : std_logic;
  signal ir20b                        : std_logic;
  signal ir21                         : std_logic;
  signal ir21b                        : std_logic;
  signal ir22                         : std_logic;
  signal ir22b                        : std_logic;
  signal ir23                         : std_logic;
  signal ir24                         : std_logic;
  signal ir25                         : std_logic;
  signal ir26                         : std_logic;
  signal ir27                         : std_logic;
  signal ir28                         : std_logic;
  signal ir29                         : std_logic;
  signal ir2                          : std_logic;
  signal ir30                         : std_logic;
  signal ir31                         : std_logic;
  signal ir32                         : std_logic;
  signal ir33                         : std_logic;
  signal ir34                         : std_logic;
  signal ir35                         : std_logic;
  signal ir36                         : std_logic;
  signal ir37                         : std_logic;
  signal ir38                         : std_logic;
  signal ir39                         : std_logic;
  signal ir3                          : std_logic;
  signal ir40                         : std_logic;
  signal ir41                         : std_logic;
  signal ir42                         : std_logic;
  signal ir43                         : std_logic;
  signal ir44                         : std_logic;
  signal ir45                         : std_logic;
  signal ir46                         : std_logic;
  signal ir47                         : std_logic;
  signal ir48                         : std_logic;
  signal ir4                          : std_logic;
  signal ir5                          : std_logic;
  signal ir6                          : std_logic;
  signal ir7                          : std_logic;
  signal ir8                          : std_logic;
  signal ir8b                         : std_logic;
  signal ir9                          : std_logic;
  signal ir9b                         : std_logic;
  signal iralu                        : std_logic;
  signal irdisp                       : std_logic;
  signal irjump                       : std_logic;
  signal iwr0                         : std_logic;
  signal iwr10                        : std_logic;
  signal iwr11                        : std_logic;
  signal iwr12                        : std_logic;
  signal iwr13                        : std_logic;
  signal iwr14                        : std_logic;
  signal iwr15                        : std_logic;
  signal iwr16                        : std_logic;
  signal iwr17                        : std_logic;
  signal iwr18                        : std_logic;
  signal iwr19                        : std_logic;
  signal iwr1                         : std_logic;
  signal iwr20                        : std_logic;
  signal iwr21                        : std_logic;
  signal iwr22                        : std_logic;
  signal iwr23                        : std_logic;
  signal iwr24                        : std_logic;
  signal iwr25                        : std_logic;
  signal iwr26                        : std_logic;
  signal iwr27                        : std_logic;
  signal iwr28                        : std_logic;
  signal iwr29                        : std_logic;
  signal iwr2                         : std_logic;
  signal iwr30                        : std_logic;
  signal iwr31                        : std_logic;
  signal iwr32                        : std_logic;
  signal iwr33                        : std_logic;
  signal iwr34                        : std_logic;
  signal iwr35                        : std_logic;
  signal iwr36                        : std_logic;
  signal iwr37                        : std_logic;
  signal iwr38                        : std_logic;
  signal iwr39                        : std_logic;
  signal iwr3                         : std_logic;
  signal iwr40                        : std_logic;
  signal iwr41                        : std_logic;
  signal iwr42                        : std_logic;
  signal iwr43                        : std_logic;
  signal iwr44                        : std_logic;
  signal iwr45                        : std_logic;
  signal iwr46                        : std_logic;
  signal iwr47                        : std_logic;
  signal iwr48                        : std_logic;
  signal iwr4                         : std_logic;
  signal iwr5                         : std_logic;
  signal iwr6                         : std_logic;
  signal iwr7                         : std_logic;
  signal iwr8                         : std_logic;
  signal iwr9                         : std_logic;
  signal iwrite                       : std_logic;
  signal iwrited                      : std_logic;
  signal iwriteda                     : std_logic;
  signal iwritedb                     : std_logic;
  signal iwritedc                     : std_logic;
  signal iwritedd                     : std_logic;
  signal iwrp1                        : std_logic;
  signal iwrp2                        : std_logic;
  signal iwrp3                        : std_logic;
  signal iwrp4                        : std_logic;
  signal jcalf                        : std_logic;
  signal jcond                        : std_logic;
  signal jfalse                       : std_logic;
  signal jret                         : std_logic;
  signal jretf                        : std_logic;
  signal l0                           : std_logic;
  signal l10                          : std_logic;
  signal l11                          : std_logic;
  signal l12                          : std_logic;
  signal l13                          : std_logic;
  signal l14                          : std_logic;
  signal l15                          : std_logic;
  signal l16                          : std_logic;
  signal l17                          : std_logic;
  signal l18                          : std_logic;
  signal l19                          : std_logic;
  signal l1                           : std_logic;
  signal l20                          : std_logic;
  signal l21                          : std_logic;
  signal l22                          : std_logic;
  signal l23                          : std_logic;
  signal l24                          : std_logic;
  signal l25                          : std_logic;
  signal l26                          : std_logic;
  signal l27                          : std_logic;
  signal l28                          : std_logic;
  signal l29                          : std_logic;
  signal l2                           : std_logic;
  signal l30                          : std_logic;
  signal l31                          : std_logic;
  signal l3                           : std_logic;
  signal l4                           : std_logic;
  signal l5                           : std_logic;
  signal l6                           : std_logic;
  signal l7                           : std_logic;
  signal l8                           : std_logic;
  signal l9                           : std_logic;
  signal lc0                          : std_logic;
  signal lc0b                         : std_logic;
  signal lc10                         : std_logic;
  signal lc11                         : std_logic;
  signal lc12                         : std_logic;
  signal lc13                         : std_logic;
  signal lc14                         : std_logic;
  signal lc15                         : std_logic;
  signal lc16                         : std_logic;
  signal lc17                         : std_logic;
  signal lc18                         : std_logic;
  signal lc19                         : std_logic;
  signal lc1                          : std_logic;
  signal lc20                         : std_logic;
  signal lc21                         : std_logic;
  signal lc22                         : std_logic;
  signal lc23                         : std_logic;
  signal lc24                         : std_logic;
  signal lc25                         : std_logic;
  signal lc2                          : std_logic;
  signal lc3                          : std_logic;
  signal lc4                          : std_logic;
  signal lc5                          : std_logic;
  signal lc6                          : std_logic;
  signal lc7                          : std_logic;
  signal lc8                          : std_logic;
  signal lc9                          : std_logic;
  signal lca0                         : std_logic;
  signal lca1                         : std_logic;
  signal lca2                         : std_logic;
  signal lca3                         : std_logic;
  signal lcdrive                      : std_logic;
  signal lcinc                        : std_logic;
  signal lcry3                        : std_logic;
  signal ldmode                       : std_logic;
  signal ldstat                       : std_logic;
  signal loadmd                       : std_logic;
  signal lparity                      : std_logic;
  signal lparl                        : std_logic;
  signal lpc0                         : std_logic;
  signal lpc10                        : std_logic;
  signal lpc11                        : std_logic;
  signal lpc12                        : std_logic;
  signal lpc13                        : std_logic;
  signal lpc1                         : std_logic;
  signal lpc2                         : std_logic;
  signal lpc3                         : std_logic;
  signal lpc4                         : std_logic;
  signal lpc5                         : std_logic;
  signal lpc6                         : std_logic;
  signal lpc7                         : std_logic;
  signal lpc8                         : std_logic;
  signal lpc9                         : std_logic;
  signal m0                           : std_logic;
  signal m10                          : std_logic;
  signal m11                          : std_logic;
  signal m12                          : std_logic;
  signal m13                          : std_logic;
  signal m14                          : std_logic;
  signal m15                          : std_logic;
  signal m16                          : std_logic;
  signal m17                          : std_logic;
  signal m18                          : std_logic;
  signal m19                          : std_logic;
  signal m1                           : std_logic;
  signal m20                          : std_logic;
  signal m21                          : std_logic;
  signal m22                          : std_logic;
  signal m23                          : std_logic;
  signal m24                          : std_logic;
  signal m25                          : std_logic;
  signal m26                          : std_logic;
  signal m27                          : std_logic;
  signal m28                          : std_logic;
  signal m29                          : std_logic;
  signal m2                           : std_logic;
  signal m30                          : std_logic;
  signal m31                          : std_logic;
  signal m31b                         : std_logic;
  signal m3                           : std_logic;
  signal m4                           : std_logic;
  signal m5                           : std_logic;
  signal m6                           : std_logic;
  signal m7                           : std_logic;
  signal m8                           : std_logic;
  signal m9                           : std_logic;
  signal machrun                      : std_logic;
  signal mapi10                       : std_logic;
  signal mapi11                       : std_logic;
  signal mapi12                       : std_logic;
  signal mapi13                       : std_logic;
  signal mapi14                       : std_logic;
  signal mapi15                       : std_logic;
  signal mapi16                       : std_logic;
  signal mapi17                       : std_logic;
  signal mapi18                       : std_logic;
  signal mapi19                       : std_logic;
  signal mapi20                       : std_logic;
  signal mapi21                       : std_logic;
  signal mapi22                       : std_logic;
  signal mapi23                       : std_logic;
  signal mapi8                        : std_logic;
  signal mapi9                        : std_logic;
  signal mapwr0d                      : std_logic;
  signal mapwr1d                      : std_logic;
  signal mbusy                        : std_logic;
  signal mclk1                        : std_logic;
  signal mclk1a                       : std_logic;
  signal mclk5                        : std_logic;
  signal mclk5a                       : std_logic;
  signal mclk7                        : std_logic;
  signal mdclk                        : std_logic;
  signal mdgetspar                    : std_logic;
  signal mdhaspar                     : std_logic;
  signal mdpar                        : std_logic;
  signal mdparerr                     : std_logic;
  signal mdpareven                    : std_logic;
  signal mdparl                       : std_logic;
  signal mdparm                       : std_logic;
  signal mdparodd                     : std_logic;
  signal mdsela                       : std_logic;
  signal mdselb                       : std_logic;
  signal mem0                         : std_logic;
  signal mem10                        : std_logic;
  signal mem11                        : std_logic;
  signal mem12                        : std_logic;
  signal mem13                        : std_logic;
  signal mem14                        : std_logic;
  signal mem15                        : std_logic;
  signal mem16                        : std_logic;
  signal mem17                        : std_logic;
  signal mem18                        : std_logic;
  signal mem19                        : std_logic;
  signal mem1                         : std_logic;
  signal mem20                        : std_logic;
  signal mem21                        : std_logic;
  signal mem22                        : std_logic;
  signal mem23                        : std_logic;
  signal mem24                        : std_logic;
  signal mem25                        : std_logic;
  signal mem26                        : std_logic;
  signal mem27                        : std_logic;
  signal mem28                        : std_logic;
  signal mem29                        : std_logic;
  signal mem2                         : std_logic;
  signal mem30                        : std_logic;
  signal mem31                        : std_logic;
  signal mem3                         : std_logic;
  signal mem4                         : std_logic;
  signal mem5                         : std_logic;
  signal mem6                         : std_logic;
  signal mem7                         : std_logic;
  signal mem8                         : std_logic;
  signal mem9                         : std_logic;
  signal memparok                     : std_logic;
  signal memprepare                   : std_logic;
  signal memrq                        : std_logic;
  signal memstart                     : std_logic;
  signal mf0                          : std_logic;
  signal mf10                         : std_logic;
  signal mf11                         : std_logic;
  signal mf12                         : std_logic;
  signal mf13                         : std_logic;
  signal mf14                         : std_logic;
  signal mf15                         : std_logic;
  signal mf16                         : std_logic;
  signal mf17                         : std_logic;
  signal mf18                         : std_logic;
  signal mf19                         : std_logic;
  signal mf1                          : std_logic;
  signal mf20                         : std_logic;
  signal mf21                         : std_logic;
  signal mf22                         : std_logic;
  signal mf23                         : std_logic;
  signal mf24                         : std_logic;
  signal mf25                         : std_logic;
  signal mf26                         : std_logic;
  signal mf27                         : std_logic;
  signal mf28                         : std_logic;
  signal mf29                         : std_logic;
  signal mf2                          : std_logic;
  signal mf30                         : std_logic;
  signal mf31                         : std_logic;
  signal mf3                          : std_logic;
  signal mf4                          : std_logic;
  signal mf5                          : std_logic;
  signal mf6                          : std_logic;
  signal mf7                          : std_logic;
  signal mf8                          : std_logic;
  signal mf9                          : std_logic;
  signal mfdrive                      : std_logic;
  signal mfenb                        : std_logic;
  signal mmem0                        : std_logic;
  signal mmem10                       : std_logic;
  signal mmem11                       : std_logic;
  signal mmem12                       : std_logic;
  signal mmem13                       : std_logic;
  signal mmem14                       : std_logic;
  signal mmem15                       : std_logic;
  signal mmem16                       : std_logic;
  signal mmem17                       : std_logic;
  signal mmem18                       : std_logic;
  signal mmem19                       : std_logic;
  signal mmem1                        : std_logic;
  signal mmem20                       : std_logic;
  signal mmem21                       : std_logic;
  signal mmem22                       : std_logic;
  signal mmem23                       : std_logic;
  signal mmem24                       : std_logic;
  signal mmem25                       : std_logic;
  signal mmem26                       : std_logic;
  signal mmem27                       : std_logic;
  signal mmem28                       : std_logic;
  signal mmem29                       : std_logic;
  signal mmem2                        : std_logic;
  signal mmem30                       : std_logic;
  signal mmem31                       : std_logic;
  signal mmem3                        : std_logic;
  signal mmem4                        : std_logic;
  signal mmem5                        : std_logic;
  signal mmem6                        : std_logic;
  signal mmem7                        : std_logic;
  signal mmem8                        : std_logic;
  signal mmem9                        : std_logic;
  signal mmemparity                   : std_logic;
  signal mmemparok                    : std_logic;
  signal mpareven                     : std_logic;
  signal mparity                      : std_logic;
  signal mparl                        : std_logic;
  signal mparm                        : std_logic;
  signal mparodd                      : std_logic;
  signal mpass                        : std_logic;
  signal mpassl                       : std_logic;
  signal msk0                         : std_logic;
  signal msk10                        : std_logic;
  signal msk11                        : std_logic;
  signal msk12                        : std_logic;
  signal msk13                        : std_logic;
  signal msk14                        : std_logic;
  signal msk15                        : std_logic;
  signal msk16                        : std_logic;
  signal msk17                        : std_logic;
  signal msk18                        : std_logic;
  signal msk19                        : std_logic;
  signal msk1                         : std_logic;
  signal msk20                        : std_logic;
  signal msk21                        : std_logic;
  signal msk22                        : std_logic;
  signal msk23                        : std_logic;
  signal msk24                        : std_logic;
  signal msk25                        : std_logic;
  signal msk26                        : std_logic;
  signal msk27                        : std_logic;
  signal msk28                        : std_logic;
  signal msk29                        : std_logic;
  signal msk2                         : std_logic;
  signal msk30                        : std_logic;
  signal msk31                        : std_logic;
  signal msk3                         : std_logic;
  signal msk4                         : std_logic;
  signal msk5                         : std_logic;
  signal msk6                         : std_logic;
  signal msk7                         : std_logic;
  signal msk8                         : std_logic;
  signal msk9                         : std_logic;
  signal mskl0                        : std_logic;
  signal mskl1                        : std_logic;
  signal mskl2                        : std_logic;
  signal mskl3                        : std_logic;
  signal mskl3cry                     : std_logic;
  signal mskl4                        : std_logic;
  signal mskr0                        : std_logic;
  signal mskr1                        : std_logic;
  signal mskr2                        : std_logic;
  signal mskr3                        : std_logic;
  signal mskr4                        : std_logic;
  signal n                            : std_logic;
  signal nc100                        : std_logic;
  signal nc101                        : std_logic;
  signal nc102                        : std_logic;
  signal nc103                        : std_logic;
  signal nc104                        : std_logic;
  signal nc105                        : std_logic;
  signal nc106                        : std_logic;
  signal nc107                        : std_logic;
  signal nc108                        : std_logic;
  signal nc109                        : std_logic;
  signal nc10                         : std_logic;
  signal nc110                        : std_logic;
  signal nc111                        : std_logic;
  signal nc112                        : std_logic;
  signal nc113                        : std_logic;
  signal nc114                        : std_logic;
  signal nc115                        : std_logic;
  signal nc116                        : std_logic;
  signal nc117                        : std_logic;
  signal nc118                        : std_logic;
  signal nc119                        : std_logic;
  signal nc11                         : std_logic;
  signal nc120                        : std_logic;
  signal nc121                        : std_logic;
  signal nc122                        : std_logic;
  signal nc123                        : std_logic;
  signal nc124                        : std_logic;
  signal nc125                        : std_logic;
  signal nc126                        : std_logic;
  signal nc127                        : std_logic;
  signal nc128                        : std_logic;
  signal nc129                        : std_logic;
  signal nc12                         : std_logic;
  signal nc130                        : std_logic;
  signal nc131                        : std_logic;
  signal nc132                        : std_logic;
  signal nc133                        : std_logic;
  signal nc134                        : std_logic;
  signal nc135                        : std_logic;
  signal nc136                        : std_logic;
  signal nc137                        : std_logic;
  signal nc138                        : std_logic;
  signal nc139                        : std_logic;
  signal nc13                         : std_logic;
  signal nc140                        : std_logic;
  signal nc141                        : std_logic;
  signal nc142                        : std_logic;
  signal nc143                        : std_logic;
  signal nc144                        : std_logic;
  signal nc145                        : std_logic;
  signal nc146                        : std_logic;
  signal nc147                        : std_logic;
  signal nc148                        : std_logic;
  signal nc149                        : std_logic;
  signal nc14                         : std_logic;
  signal nc150                        : std_logic;
  signal nc151                        : std_logic;
  signal nc152                        : std_logic;
  signal nc153                        : std_logic;
  signal nc154                        : std_logic;
  signal nc155                        : std_logic;
  signal nc156                        : std_logic;
  signal nc157                        : std_logic;
  signal nc158                        : std_logic;
  signal nc159                        : std_logic;
  signal nc15                         : std_logic;
  signal nc160                        : std_logic;
  signal nc161                        : std_logic;
  signal nc162                        : std_logic;
  signal nc163                        : std_logic;
  signal nc164                        : std_logic;
  signal nc165                        : std_logic;
  signal nc166                        : std_logic;
  signal nc167                        : std_logic;
  signal nc168                        : std_logic;
  signal nc169                        : std_logic;
  signal nc16                         : std_logic;
  signal nc170                        : std_logic;
  signal nc171                        : std_logic;
  signal nc172                        : std_logic;
  signal nc173                        : std_logic;
  signal nc174                        : std_logic;
  signal nc175                        : std_logic;
  signal nc176                        : std_logic;
  signal nc177                        : std_logic;
  signal nc178                        : std_logic;
  signal nc179                        : std_logic;
  signal nc17                         : std_logic;
  signal nc180                        : std_logic;
  signal nc181                        : std_logic;
  signal nc182                        : std_logic;
  signal nc183                        : std_logic;
  signal nc184                        : std_logic;
  signal nc185                        : std_logic;
  signal nc186                        : std_logic;
  signal nc187                        : std_logic;
  signal nc188                        : std_logic;
  signal nc189                        : std_logic;
  signal nc18                         : std_logic;
  signal nc190                        : std_logic;
  signal nc191                        : std_logic;
  signal nc192                        : std_logic;
  signal nc193                        : std_logic;
  signal nc194                        : std_logic;
  signal nc195                        : std_logic;
  signal nc196                        : std_logic;
  signal nc197                        : std_logic;
  signal nc198                        : std_logic;
  signal nc199                        : std_logic;
  signal nc19                         : std_logic;
  signal nc1                          : std_logic;
  signal nc200                        : std_logic;
  signal nc201                        : std_logic;
  signal nc202                        : std_logic;
  signal nc203                        : std_logic;
  signal nc204                        : std_logic;
  signal nc205                        : std_logic;
  signal nc206                        : std_logic;
  signal nc207                        : std_logic;
  signal nc208                        : std_logic;
  signal nc209                        : std_logic;
  signal nc20                         : std_logic;
  signal nc210                        : std_logic;
  signal nc211                        : std_logic;
  signal nc212                        : std_logic;
  signal nc213                        : std_logic;
  signal nc214                        : std_logic;
  signal nc215                        : std_logic;
  signal nc216                        : std_logic;
  signal nc217                        : std_logic;
  signal nc218                        : std_logic;
  signal nc219                        : std_logic;
  signal nc21                         : std_logic;
  signal nc220                        : std_logic;
  signal nc221                        : std_logic;
  signal nc222                        : std_logic;
  signal nc223                        : std_logic;
  signal nc224                        : std_logic;
  signal nc225                        : std_logic;
  signal nc226                        : std_logic;
  signal nc227                        : std_logic;
  signal nc228                        : std_logic;
  signal nc229                        : std_logic;
  signal nc22                         : std_logic;
  signal nc230                        : std_logic;
  signal nc231                        : std_logic;
  signal nc232                        : std_logic;
  signal nc233                        : std_logic;
  signal nc234                        : std_logic;
  signal nc235                        : std_logic;
  signal nc236                        : std_logic;
  signal nc237                        : std_logic;
  signal nc238                        : std_logic;
  signal nc239                        : std_logic;
  signal nc23                         : std_logic;
  signal nc240                        : std_logic;
  signal nc241                        : std_logic;
  signal nc242                        : std_logic;
  signal nc243                        : std_logic;
  signal nc244                        : std_logic;
  signal nc245                        : std_logic;
  signal nc246                        : std_logic;
  signal nc247                        : std_logic;
  signal nc248                        : std_logic;
  signal nc249                        : std_logic;
  signal nc24                         : std_logic;
  signal nc250                        : std_logic;
  signal nc251                        : std_logic;
  signal nc252                        : std_logic;
  signal nc253                        : std_logic;
  signal nc254                        : std_logic;
  signal nc255                        : std_logic;
  signal nc256                        : std_logic;
  signal nc257                        : std_logic;
  signal nc258                        : std_logic;
  signal nc259                        : std_logic;
  signal nc25                         : std_logic;
  signal nc260                        : std_logic;
  signal nc261                        : std_logic;
  signal nc262                        : std_logic;
  signal nc263                        : std_logic;
  signal nc264                        : std_logic;
  signal nc265                        : std_logic;
  signal nc266                        : std_logic;
  signal nc267                        : std_logic;
  signal nc268                        : std_logic;
  signal nc269                        : std_logic;
  signal nc26                         : std_logic;
  signal nc270                        : std_logic;
  signal nc271                        : std_logic;
  signal nc272                        : std_logic;
  signal nc273                        : std_logic;
  signal nc274                        : std_logic;
  signal nc275                        : std_logic;
  signal nc276                        : std_logic;
  signal nc277                        : std_logic;
  signal nc278                        : std_logic;
  signal nc279                        : std_logic;
  signal nc27                         : std_logic;
  signal nc280                        : std_logic;
  signal nc281                        : std_logic;
  signal nc282                        : std_logic;
  signal nc283                        : std_logic;
  signal nc284                        : std_logic;
  signal nc285                        : std_logic;
  signal nc286                        : std_logic;
  signal nc287                        : std_logic;
  signal nc288                        : std_logic;
  signal nc289                        : std_logic;
  signal nc28                         : std_logic;
  signal nc290                        : std_logic;
  signal nc291                        : std_logic;
  signal nc292                        : std_logic;
  signal nc293                        : std_logic;
  signal nc294                        : std_logic;
  signal nc295                        : std_logic;
  signal nc296                        : std_logic;
  signal nc297                        : std_logic;
  signal nc298                        : std_logic;
  signal nc299                        : std_logic;
  signal nc29                         : std_logic;
  signal nc2                          : std_logic;
  signal nc300                        : std_logic;
  signal nc301                        : std_logic;
  signal nc302                        : std_logic;
  signal nc303                        : std_logic;
  signal nc304                        : std_logic;
  signal nc305                        : std_logic;
  signal nc306                        : std_logic;
  signal nc307                        : std_logic;
  signal nc308                        : std_logic;
  signal nc309                        : std_logic;
  signal nc30                         : std_logic;
  signal nc310                        : std_logic;
  signal nc311                        : std_logic;
  signal nc312                        : std_logic;
  signal nc313                        : std_logic;
  signal nc314                        : std_logic;
  signal nc315                        : std_logic;
  signal nc316                        : std_logic;
  signal nc317                        : std_logic;
  signal nc318                        : std_logic;
  signal nc319                        : std_logic;
  signal nc31                         : std_logic;
  signal nc320                        : std_logic;
  signal nc321                        : std_logic;
  signal nc322                        : std_logic;
  signal nc323                        : std_logic;
  signal nc324                        : std_logic;
  signal nc325                        : std_logic;
  signal nc326                        : std_logic;
  signal nc327                        : std_logic;
  signal nc328                        : std_logic;
  signal nc329                        : std_logic;
  signal nc32                         : std_logic;
  signal nc330                        : std_logic;
  signal nc331                        : std_logic;
  signal nc332                        : std_logic;
  signal nc333                        : std_logic;
  signal nc334                        : std_logic;
  signal nc335                        : std_logic;
  signal nc336                        : std_logic;
  signal nc337                        : std_logic;
  signal nc338                        : std_logic;
  signal nc339                        : std_logic;
  signal nc33                         : std_logic;
  signal nc340                        : std_logic;
  signal nc341                        : std_logic;
  signal nc342                        : std_logic;
  signal nc343                        : std_logic;
  signal nc344                        : std_logic;
  signal nc345                        : std_logic;
  signal nc346                        : std_logic;
  signal nc347                        : std_logic;
  signal nc348                        : std_logic;
  signal nc349                        : std_logic;
  signal nc34                         : std_logic;
  signal nc350                        : std_logic;
  signal nc351                        : std_logic;
  signal nc352                        : std_logic;
  signal nc353                        : std_logic;
  signal nc354                        : std_logic;
  signal nc355                        : std_logic;
  signal nc356                        : std_logic;
  signal nc357                        : std_logic;
  signal nc358                        : std_logic;
  signal nc359                        : std_logic;
  signal nc35                         : std_logic;
  signal nc360                        : std_logic;
  signal nc361                        : std_logic;
  signal nc362                        : std_logic;
  signal nc363                        : std_logic;
  signal nc364                        : std_logic;
  signal nc365                        : std_logic;
  signal nc366                        : std_logic;
  signal nc367                        : std_logic;
  signal nc368                        : std_logic;
  signal nc369                        : std_logic;
  signal nc36                         : std_logic;
  signal nc370                        : std_logic;
  signal nc371                        : std_logic;
  signal nc372                        : std_logic;
  signal nc373                        : std_logic;
  signal nc374                        : std_logic;
  signal nc375                        : std_logic;
  signal nc376                        : std_logic;
  signal nc377                        : std_logic;
  signal nc378                        : std_logic;
  signal nc379                        : std_logic;
  signal nc37                         : std_logic;
  signal nc380                        : std_logic;
  signal nc381                        : std_logic;
  signal nc382                        : std_logic;
  signal nc383                        : std_logic;
  signal nc384                        : std_logic;
  signal nc385                        : std_logic;
  signal nc386                        : std_logic;
  signal nc387                        : std_logic;
  signal nc388                        : std_logic;
  signal nc389                        : std_logic;
  signal nc38                         : std_logic;
  signal nc390                        : std_logic;
  signal nc391                        : std_logic;
  signal nc392                        : std_logic;
  signal nc393                        : std_logic;
  signal nc394                        : std_logic;
  signal nc395                        : std_logic;
  signal nc396                        : std_logic;
  signal nc397                        : std_logic;
  signal nc398                        : std_logic;
  signal nc399                        : std_logic;
  signal nc39                         : std_logic;
  signal nc3                          : std_logic;
  signal nc400                        : std_logic;
  signal nc401                        : std_logic;
  signal nc402                        : std_logic;
  signal nc403                        : std_logic;
  signal nc404                        : std_logic;
  signal nc405                        : std_logic;
  signal nc406                        : std_logic;
  signal nc407                        : std_logic;
  signal nc408                        : std_logic;
  signal nc409                        : std_logic;
  signal nc40                         : std_logic;
  signal nc410                        : std_logic;
  signal nc411                        : std_logic;
  signal nc412                        : std_logic;
  signal nc413                        : std_logic;
  signal nc414                        : std_logic;
  signal nc415                        : std_logic;
  signal nc416                        : std_logic;
  signal nc417                        : std_logic;
  signal nc418                        : std_logic;
  signal nc419                        : std_logic;
  signal nc41                         : std_logic;
  signal nc420                        : std_logic;
  signal nc421                        : std_logic;
  signal nc422                        : std_logic;
  signal nc423                        : std_logic;
  signal nc424                        : std_logic;
  signal nc425                        : std_logic;
  signal nc426                        : std_logic;
  signal nc427                        : std_logic;
  signal nc428                        : std_logic;
  signal nc429                        : std_logic;
  signal nc42                         : std_logic;
  signal nc430                        : std_logic;
  signal nc431                        : std_logic;
  signal nc432                        : std_logic;
  signal nc433                        : std_logic;
  signal nc434                        : std_logic;
  signal nc435                        : std_logic;
  signal nc436                        : std_logic;
  signal nc437                        : std_logic;
  signal nc438                        : std_logic;
  signal nc439                        : std_logic;
  signal nc43                         : std_logic;
  signal nc440                        : std_logic;
  signal nc441                        : std_logic;
  signal nc442                        : std_logic;
  signal nc443                        : std_logic;
  signal nc444                        : std_logic;
  signal nc445                        : std_logic;
  signal nc446                        : std_logic;
  signal nc447                        : std_logic;
  signal nc448                        : std_logic;
  signal nc449                        : std_logic;
  signal nc44                         : std_logic;
  signal nc450                        : std_logic;
  signal nc451                        : std_logic;
  signal nc452                        : std_logic;
  signal nc453                        : std_logic;
  signal nc454                        : std_logic;
  signal nc455                        : std_logic;
  signal nc456                        : std_logic;
  signal nc457                        : std_logic;
  signal nc458                        : std_logic;
  signal nc459                        : std_logic;
  signal nc45                         : std_logic;
  signal nc460                        : std_logic;
  signal nc461                        : std_logic;
  signal nc462                        : std_logic;
  signal nc463                        : std_logic;
  signal nc464                        : std_logic;
  signal nc465                        : std_logic;
  signal nc466                        : std_logic;
  signal nc467                        : std_logic;
  signal nc468                        : std_logic;
  signal nc469                        : std_logic;
  signal nc46                         : std_logic;
  signal nc470                        : std_logic;
  signal nc471                        : std_logic;
  signal nc472                        : std_logic;
  signal nc473                        : std_logic;
  signal nc474                        : std_logic;
  signal nc475                        : std_logic;
  signal nc476                        : std_logic;
  signal nc477                        : std_logic;
  signal nc478                        : std_logic;
  signal nc479                        : std_logic;
  signal nc47                         : std_logic;
  signal nc480                        : std_logic;
  signal nc481                        : std_logic;
  signal nc482                        : std_logic;
  signal nc483                        : std_logic;
  signal nc484                        : std_logic;
  signal nc485                        : std_logic;
  signal nc486                        : std_logic;
  signal nc487                        : std_logic;
  signal nc488                        : std_logic;
  signal nc489                        : std_logic;
  signal nc48                         : std_logic;
  signal nc490                        : std_logic;
  signal nc491                        : std_logic;
  signal nc492                        : std_logic;
  signal nc493                        : std_logic;
  signal nc494                        : std_logic;
  signal nc49                         : std_logic;
  signal nc4                          : std_logic;
  signal nc50                         : std_logic;
  signal nc51                         : std_logic;
  signal nc52                         : std_logic;
  signal nc53                         : std_logic;
  signal nc54                         : std_logic;
  signal nc55                         : std_logic;
  signal nc56                         : std_logic;
  signal nc57                         : std_logic;
  signal nc58                         : std_logic;
  signal nc59                         : std_logic;
  signal nc5                          : std_logic;
  signal nc60                         : std_logic;
  signal nc61                         : std_logic;
  signal nc62                         : std_logic;
  signal nc63                         : std_logic;
  signal nc64                         : std_logic;
  signal nc65                         : std_logic;
  signal nc66                         : std_logic;
  signal nc67                         : std_logic;
  signal nc68                         : std_logic;
  signal nc69                         : std_logic;
  signal nc6                          : std_logic;
  signal nc70                         : std_logic;
  signal nc71                         : std_logic;
  signal nc72                         : std_logic;
  signal nc73                         : std_logic;
  signal nc74                         : std_logic;
  signal nc75                         : std_logic;
  signal nc76                         : std_logic;
  signal nc77                         : std_logic;
  signal nc78                         : std_logic;
  signal nc79                         : std_logic;
  signal nc7                          : std_logic;
  signal nc80                         : std_logic;
  signal nc81                         : std_logic;
  signal nc82                         : std_logic;
  signal nc83                         : std_logic;
  signal nc84                         : std_logic;
  signal nc85                         : std_logic;
  signal nc86                         : std_logic;
  signal nc87                         : std_logic;
  signal nc88                         : std_logic;
  signal nc89                         : std_logic;
  signal nc8                          : std_logic;
  signal nc90                         : std_logic;
  signal nc91                         : std_logic;
  signal nc92                         : std_logic;
  signal nc93                         : std_logic;
  signal nc94                         : std_logic;
  signal nc95                         : std_logic;
  signal nc96                         : std_logic;
  signal nc97                         : std_logic;
  signal nc98                         : std_logic;
  signal nc99                         : std_logic;
  signal nc9                          : std_logic;
  signal needfetch                    : std_logic;
  signal newlc                        : std_logic;
  signal nop11                        : std_logic;
  signal nop                          : std_logic;
  signal nopa                         : std_logic;
  signal npc0                         : std_logic;
  signal npc10                        : std_logic;
  signal npc11                        : std_logic;
  signal npc12                        : std_logic;
  signal npc13                        : std_logic;
  signal npc1                         : std_logic;
  signal npc2                         : std_logic;
  signal npc3                         : std_logic;
  signal npc4                         : std_logic;
  signal npc5                         : std_logic;
  signal npc6                         : std_logic;
  signal npc7                         : std_logic;
  signal npc8                         : std_logic;
  signal npc9                         : std_logic;
  signal ob0                          : std_logic;
  signal ob10                         : std_logic;
  signal ob11                         : std_logic;
  signal ob12                         : std_logic;
  signal ob13                         : std_logic;
  signal ob14                         : std_logic;
  signal ob15                         : std_logic;
  signal ob16                         : std_logic;
  signal ob17                         : std_logic;
  signal ob18                         : std_logic;
  signal ob19                         : std_logic;
  signal ob1                          : std_logic;
  signal ob20                         : std_logic;
  signal ob21                         : std_logic;
  signal ob22                         : std_logic;
  signal ob23                         : std_logic;
  signal ob24                         : std_logic;
  signal ob25                         : std_logic;
  signal ob26                         : std_logic;
  signal ob27                         : std_logic;
  signal ob28                         : std_logic;
  signal ob29                         : std_logic;
  signal ob2                          : std_logic;
  signal ob30                         : std_logic;
  signal ob31                         : std_logic;
  signal ob3                          : std_logic;
  signal ob4                          : std_logic;
  signal ob5                          : std_logic;
  signal ob6                          : std_logic;
  signal ob7                          : std_logic;
  signal ob8                          : std_logic;
  signal ob9                          : std_logic;
  signal opc0                         : std_logic;
  signal opc10                        : std_logic;
  signal opc11                        : std_logic;
  signal opc12                        : std_logic;
  signal opc13                        : std_logic;
  signal opc1                         : std_logic;
  signal opc2                         : std_logic;
  signal opc3                         : std_logic;
  signal opc4                         : std_logic;
  signal opc5                         : std_logic;
  signal opc6                         : std_logic;
  signal opc7                         : std_logic;
  signal opc8                         : std_logic;
  signal opc9                         : std_logic;
  signal opcclk                       : std_logic;
  signal opcclka                      : std_logic;
  signal opcclkb                      : std_logic;
  signal opcclkc                      : std_logic;
  signal opcinh                       : std_logic;
  signal opcinha                      : std_logic;
  signal opcinhb                      : std_logic;
  signal osel0a                       : std_logic;
  signal osel0b                       : std_logic;
  signal osel1a                       : std_logic;
  signal osel1b                       : std_logic;
  signal pc0                          : std_logic;
  signal pc0a                         : std_logic;
  signal pc0b                         : std_logic;
  signal pc0c                         : std_logic;
  signal pc0d                         : std_logic;
  signal pc0e                         : std_logic;
  signal pc0f                         : std_logic;
  signal pc0g                         : std_logic;
  signal pc0h                         : std_logic;
  signal pc0i                         : std_logic;
  signal pc0j                         : std_logic;
  signal pc0k                         : std_logic;
  signal pc0l                         : std_logic;
  signal pc0m                         : std_logic;
  signal pc0n                         : std_logic;
  signal pc0o                         : std_logic;
  signal pc0p                         : std_logic;
  signal pc10                         : std_logic;
  signal pc10a                        : std_logic;
  signal pc10b                        : std_logic;
  signal pc10c                        : std_logic;
  signal pc10d                        : std_logic;
  signal pc10e                        : std_logic;
  signal pc10f                        : std_logic;
  signal pc10g                        : std_logic;
  signal pc10h                        : std_logic;
  signal pc10i                        : std_logic;
  signal pc10j                        : std_logic;
  signal pc10k                        : std_logic;
  signal pc10l                        : std_logic;
  signal pc10m                        : std_logic;
  signal pc10n                        : std_logic;
  signal pc10o                        : std_logic;
  signal pc10p                        : std_logic;
  signal pc11                         : std_logic;
  signal pc11a                        : std_logic;
  signal pc11b                        : std_logic;
  signal pc11c                        : std_logic;
  signal pc11d                        : std_logic;
  signal pc11e                        : std_logic;
  signal pc11f                        : std_logic;
  signal pc11g                        : std_logic;
  signal pc11h                        : std_logic;
  signal pc11i                        : std_logic;
  signal pc11j                        : std_logic;
  signal pc11k                        : std_logic;
  signal pc11l                        : std_logic;
  signal pc11m                        : std_logic;
  signal pc11n                        : std_logic;
  signal pc11o                        : std_logic;
  signal pc11p                        : std_logic;
  signal pc12                         : std_logic;
  signal pc12b                        : std_logic;
  signal pc13                         : std_logic;
  signal pc13b                        : std_logic;
  signal pc1                          : std_logic;
  signal pc1a                         : std_logic;
  signal pc1b                         : std_logic;
  signal pc1c                         : std_logic;
  signal pc1d                         : std_logic;
  signal pc1e                         : std_logic;
  signal pc1f                         : std_logic;
  signal pc1g                         : std_logic;
  signal pc1h                         : std_logic;
  signal pc1i                         : std_logic;
  signal pc1j                         : std_logic;
  signal pc1k                         : std_logic;
  signal pc1l                         : std_logic;
  signal pc1m                         : std_logic;
  signal pc1n                         : std_logic;
  signal pc1o                         : std_logic;
  signal pc1p                         : std_logic;
  signal pc2                          : std_logic;
  signal pc2a                         : std_logic;
  signal pc2b                         : std_logic;
  signal pc2c                         : std_logic;
  signal pc2d                         : std_logic;
  signal pc2e                         : std_logic;
  signal pc2f                         : std_logic;
  signal pc2g                         : std_logic;
  signal pc2h                         : std_logic;
  signal pc2i                         : std_logic;
  signal pc2j                         : std_logic;
  signal pc2k                         : std_logic;
  signal pc2l                         : std_logic;
  signal pc2m                         : std_logic;
  signal pc2n                         : std_logic;
  signal pc2o                         : std_logic;
  signal pc2p                         : std_logic;
  signal pc3                          : std_logic;
  signal pc3a                         : std_logic;
  signal pc3b                         : std_logic;
  signal pc3c                         : std_logic;
  signal pc3d                         : std_logic;
  signal pc3e                         : std_logic;
  signal pc3f                         : std_logic;
  signal pc3g                         : std_logic;
  signal pc3h                         : std_logic;
  signal pc3i                         : std_logic;
  signal pc3j                         : std_logic;
  signal pc3k                         : std_logic;
  signal pc3l                         : std_logic;
  signal pc3m                         : std_logic;
  signal pc3n                         : std_logic;
  signal pc3o                         : std_logic;
  signal pc3p                         : std_logic;
  signal pc4                          : std_logic;
  signal pc4a                         : std_logic;
  signal pc4b                         : std_logic;
  signal pc4c                         : std_logic;
  signal pc4d                         : std_logic;
  signal pc4e                         : std_logic;
  signal pc4f                         : std_logic;
  signal pc4g                         : std_logic;
  signal pc4h                         : std_logic;
  signal pc4i                         : std_logic;
  signal pc4j                         : std_logic;
  signal pc4k                         : std_logic;
  signal pc4l                         : std_logic;
  signal pc4m                         : std_logic;
  signal pc4n                         : std_logic;
  signal pc4o                         : std_logic;
  signal pc4p                         : std_logic;
  signal pc5                          : std_logic;
  signal pc5a                         : std_logic;
  signal pc5b                         : std_logic;
  signal pc5c                         : std_logic;
  signal pc5d                         : std_logic;
  signal pc5e                         : std_logic;
  signal pc5f                         : std_logic;
  signal pc5g                         : std_logic;
  signal pc5h                         : std_logic;
  signal pc5i                         : std_logic;
  signal pc5j                         : std_logic;
  signal pc5k                         : std_logic;
  signal pc5l                         : std_logic;
  signal pc5m                         : std_logic;
  signal pc5n                         : std_logic;
  signal pc5o                         : std_logic;
  signal pc5p                         : std_logic;
  signal pc6                          : std_logic;
  signal pc6a                         : std_logic;
  signal pc6b                         : std_logic;
  signal pc6c                         : std_logic;
  signal pc6d                         : std_logic;
  signal pc6e                         : std_logic;
  signal pc6f                         : std_logic;
  signal pc6g                         : std_logic;
  signal pc6h                         : std_logic;
  signal pc6i                         : std_logic;
  signal pc6j                         : std_logic;
  signal pc6k                         : std_logic;
  signal pc6l                         : std_logic;
  signal pc6m                         : std_logic;
  signal pc6n                         : std_logic;
  signal pc6o                         : std_logic;
  signal pc6p                         : std_logic;
  signal pc7                          : std_logic;
  signal pc7a                         : std_logic;
  signal pc7b                         : std_logic;
  signal pc7c                         : std_logic;
  signal pc7d                         : std_logic;
  signal pc7e                         : std_logic;
  signal pc7f                         : std_logic;
  signal pc7g                         : std_logic;
  signal pc7h                         : std_logic;
  signal pc7i                         : std_logic;
  signal pc7j                         : std_logic;
  signal pc7k                         : std_logic;
  signal pc7l                         : std_logic;
  signal pc7m                         : std_logic;
  signal pc7n                         : std_logic;
  signal pc7o                         : std_logic;
  signal pc7p                         : std_logic;
  signal pc8                          : std_logic;
  signal pc8a                         : std_logic;
  signal pc8b                         : std_logic;
  signal pc8c                         : std_logic;
  signal pc8d                         : std_logic;
  signal pc8e                         : std_logic;
  signal pc8f                         : std_logic;
  signal pc8g                         : std_logic;
  signal pc8h                         : std_logic;
  signal pc8i                         : std_logic;
  signal pc8j                         : std_logic;
  signal pc8k                         : std_logic;
  signal pc8l                         : std_logic;
  signal pc8m                         : std_logic;
  signal pc8n                         : std_logic;
  signal pc8o                         : std_logic;
  signal pc8p                         : std_logic;
  signal pc9                          : std_logic;
  signal pc9a                         : std_logic;
  signal pc9b                         : std_logic;
  signal pc9c                         : std_logic;
  signal pc9d                         : std_logic;
  signal pc9e                         : std_logic;
  signal pc9f                         : std_logic;
  signal pc9g                         : std_logic;
  signal pc9h                         : std_logic;
  signal pc9i                         : std_logic;
  signal pc9j                         : std_logic;
  signal pc9k                         : std_logic;
  signal pc9l                         : std_logic;
  signal pc9m                         : std_logic;
  signal pc9n                         : std_logic;
  signal pc9o                         : std_logic;
  signal pc9p                         : std_logic;
  signal pccry11                      : std_logic;
  signal pccry3                       : std_logic;
  signal pccry7                       : std_logic;
  signal pcs0                         : std_logic;
  signal pcs1                         : std_logic;
  signal pdl0                         : std_logic;
  signal pdl10                        : std_logic;
  signal pdl11                        : std_logic;
  signal pdl12                        : std_logic;
  signal pdl13                        : std_logic;
  signal pdl14                        : std_logic;
  signal pdl15                        : std_logic;
  signal pdl16                        : std_logic;
  signal pdl17                        : std_logic;
  signal pdl18                        : std_logic;
  signal pdl19                        : std_logic;
  signal pdl1                         : std_logic;
  signal pdl20                        : std_logic;
  signal pdl21                        : std_logic;
  signal pdl22                        : std_logic;
  signal pdl23                        : std_logic;
  signal pdl24                        : std_logic;
  signal pdl25                        : std_logic;
  signal pdl26                        : std_logic;
  signal pdl27                        : std_logic;
  signal pdl28                        : std_logic;
  signal pdl29                        : std_logic;
  signal pdl2                         : std_logic;
  signal pdl30                        : std_logic;
  signal pdl31                        : std_logic;
  signal pdl3                         : std_logic;
  signal pdl4                         : std_logic;
  signal pdl5                         : std_logic;
  signal pdl6                         : std_logic;
  signal pdl7                         : std_logic;
  signal pdl8                         : std_logic;
  signal pdl9                         : std_logic;
  signal pdlenb                       : std_logic;
  signal pdlidx0                      : std_logic;
  signal pdlidx1                      : std_logic;
  signal pdlidx2                      : std_logic;
  signal pdlidx3                      : std_logic;
  signal pdlidx4                      : std_logic;
  signal pdlidx5                      : std_logic;
  signal pdlidx6                      : std_logic;
  signal pdlidx7                      : std_logic;
  signal pdlidx8                      : std_logic;
  signal pdlidx9                      : std_logic;
  signal pdlparity                    : std_logic;
  signal pdlparok                     : std_logic;
  signal pdlptr0                      : std_logic;
  signal pdlptr1                      : std_logic;
  signal pdlptr2                      : std_logic;
  signal pdlptr3                      : std_logic;
  signal pdlptr4                      : std_logic;
  signal pdlptr5                      : std_logic;
  signal pdlptr6                      : std_logic;
  signal pdlptr7                      : std_logic;
  signal pdlptr8                      : std_logic;
  signal pdlptr9                      : std_logic;
  signal pdlwrite                     : std_logic;
  signal pdlwrited                    : std_logic;
  signal pidrive                      : std_logic;
  signal popj                         : std_logic;
  signal promdisable                  : std_logic;
  signal promdisabled                 : std_logic;
  signal promenable                   : std_logic;
  signal pwidx                        : std_logic;
  signal q0                           : std_logic;
  signal q10                          : std_logic;
  signal q11                          : std_logic;
  signal q12                          : std_logic;
  signal q13                          : std_logic;
  signal q14                          : std_logic;
  signal q15                          : std_logic;
  signal q16                          : std_logic;
  signal q17                          : std_logic;
  signal q18                          : std_logic;
  signal q19                          : std_logic;
  signal q1                           : std_logic;
  signal q20                          : std_logic;
  signal q21                          : std_logic;
  signal q22                          : std_logic;
  signal q23                          : std_logic;
  signal q24                          : std_logic;
  signal q25                          : std_logic;
  signal q26                          : std_logic;
  signal q27                          : std_logic;
  signal q28                          : std_logic;
  signal q29                          : std_logic;
  signal q2                           : std_logic;
  signal q30                          : std_logic;
  signal q31                          : std_logic;
  signal q3                           : std_logic;
  signal q4                           : std_logic;
  signal q5                           : std_logic;
  signal q6                           : std_logic;
  signal q7                           : std_logic;
  signal q8                           : std_logic;
  signal q9                           : std_logic;
  signal qdrive                       : std_logic;
  signal qs0                          : std_logic;
  signal qs1                          : std_logic;
  signal r0                           : std_logic;
  signal r10                          : std_logic;
  signal r11                          : std_logic;
  signal r12                          : std_logic;
  signal r13                          : std_logic;
  signal r14                          : std_logic;
  signal r15                          : std_logic;
  signal r16                          : std_logic;
  signal r17                          : std_logic;
  signal r18                          : std_logic;
  signal r19                          : std_logic;
  signal r1                           : std_logic;
  signal r20                          : std_logic;
  signal r21                          : std_logic;
  signal r22                          : std_logic;
  signal r23                          : std_logic;
  signal r24                          : std_logic;
  signal r25                          : std_logic;
  signal r26                          : std_logic;
  signal r27                          : std_logic;
  signal r28                          : std_logic;
  signal r29                          : std_logic;
  signal r2                           : std_logic;
  signal r30                          : std_logic;
  signal r31                          : std_logic;
  signal r3                           : std_logic;
  signal r4                           : std_logic;
  signal r5                           : std_logic;
  signal r6                           : std_logic;
  signal r7                           : std_logic;
  signal r8                           : std_logic;
  signal r9                           : std_logic;
  signal ramdisable                   : std_logic;
  signal rdcyc                        : std_logic;
  signal reset                        : std_logic;
  signal reta0                        : std_logic;
  signal reta10                       : std_logic;
  signal reta11                       : std_logic;
  signal reta12                       : std_logic;
  signal reta13                       : std_logic;
  signal reta1                        : std_logic;
  signal reta2                        : std_logic;
  signal reta3                        : std_logic;
  signal reta4                        : std_logic;
  signal reta5                        : std_logic;
  signal reta6                        : std_logic;
  signal reta7                        : std_logic;
  signal reta8                        : std_logic;
  signal reta9                        : std_logic;
  signal run                          : std_logic;
  signal s0                           : std_logic;
  signal s1                           : std_logic;
  signal s2a                          : std_logic;
  signal s2b                          : std_logic;
  signal s3a                          : std_logic;
  signal s3b                          : std_logic;
  signal s4                           : std_logic;
  signal sa0                          : std_logic;
  signal sa10                         : std_logic;
  signal sa11                         : std_logic;
  signal sa12                         : std_logic;
  signal sa13                         : std_logic;
  signal sa14                         : std_logic;
  signal sa15                         : std_logic;
  signal sa16                         : std_logic;
  signal sa17                         : std_logic;
  signal sa18                         : std_logic;
  signal sa19                         : std_logic;
  signal sa1                          : std_logic;
  signal sa20                         : std_logic;
  signal sa21                         : std_logic;
  signal sa22                         : std_logic;
  signal sa23                         : std_logic;
  signal sa24                         : std_logic;
  signal sa25                         : std_logic;
  signal sa26                         : std_logic;
  signal sa27                         : std_logic;
  signal sa28                         : std_logic;
  signal sa29                         : std_logic;
  signal sa2                          : std_logic;
  signal sa30                         : std_logic;
  signal sa31                         : std_logic;
  signal sa3                          : std_logic;
  signal sa4                          : std_logic;
  signal sa5                          : std_logic;
  signal sa6                          : std_logic;
  signal sa7                          : std_logic;
  signal sa8                          : std_logic;
  signal sa9                          : std_logic;
  signal sint                         : std_logic;
  signal sintr                        : std_logic;
  signal spc0                         : std_logic;
  signal spc10                        : std_logic;
  signal spc11                        : std_logic;
  signal spc12                        : std_logic;
  signal spc13                        : std_logic;
  signal spc14                        : std_logic;
  signal spc15                        : std_logic;
  signal spc16                        : std_logic;
  signal spc17                        : std_logic;
  signal spc18                        : std_logic;
  signal spc1                         : std_logic;
  signal spc1a                        : std_logic;
  signal spc2                         : std_logic;
  signal spc3                         : std_logic;
  signal spc4                         : std_logic;
  signal spc5                         : std_logic;
  signal spc6                         : std_logic;
  signal spc7                         : std_logic;
  signal spc8                         : std_logic;
  signal spc9                         : std_logic;
  signal spcdrive                     : std_logic;
  signal spcenb                       : std_logic;
  signal spcmung                      : std_logic;
  signal spco0                        : std_logic;
  signal spco10                       : std_logic;
  signal spco11                       : std_logic;
  signal spco12                       : std_logic;
  signal spco13                       : std_logic;
  signal spco14                       : std_logic;
  signal spco15                       : std_logic;
  signal spco16                       : std_logic;
  signal spco17                       : std_logic;
  signal spco18                       : std_logic;
  signal spco1                        : std_logic;
  signal spco2                        : std_logic;
  signal spco3                        : std_logic;
  signal spco4                        : std_logic;
  signal spco5                        : std_logic;
  signal spco6                        : std_logic;
  signal spco7                        : std_logic;
  signal spco8                        : std_logic;
  signal spco9                        : std_logic;
  signal spcopar                      : std_logic;
  signal spcpar                       : std_logic;
  signal spcparh                      : std_logic;
  signal spcparok                     : std_logic;
  signal spcptr0                      : std_logic;
  signal spcptr1                      : std_logic;
  signal spcptr2                      : std_logic;
  signal spcptr3                      : std_logic;
  signal spcptr4                      : std_logic;
  signal spcw0                        : std_logic;
  signal spcw10                       : std_logic;
  signal spcw11                       : std_logic;
  signal spcw12                       : std_logic;
  signal spcw13                       : std_logic;
  signal spcw14                       : std_logic;
  signal spcw15                       : std_logic;
  signal spcw16                       : std_logic;
  signal spcw17                       : std_logic;
  signal spcw18                       : std_logic;
  signal spcw1                        : std_logic;
  signal spcw2                        : std_logic;
  signal spcw3                        : std_logic;
  signal spcw4                        : std_logic;
  signal spcw5                        : std_logic;
  signal spcw6                        : std_logic;
  signal spcw7                        : std_logic;
  signal spcw8                        : std_logic;
  signal spcw9                        : std_logic;
  signal spcwpar                      : std_logic;
  signal spcwparh                     : std_logic;
  signal spcwpass                     : std_logic;
  signal speed0                       : std_logic;
  signal speed0a                      : std_logic;
  signal speed1                       : std_logic;
  signal speed1a                      : std_logic;
  signal speedclk                     : std_logic;
  signal spush                        : std_logic;
  signal spushd                       : std_logic;
  signal spy0                         : std_logic;
  signal spy10                        : std_logic;
  signal spy11                        : std_logic;
  signal spy12                        : std_logic;
  signal spy13                        : std_logic;
  signal spy14                        : std_logic;
  signal spy15                        : std_logic;
  signal spy1                         : std_logic;
  signal spy2                         : std_logic;
  signal spy3                         : std_logic;
  signal spy4                         : std_logic;
  signal spy5                         : std_logic;
  signal spy6                         : std_logic;
  signal spy7                         : std_logic;
  signal spy8                         : std_logic;
  signal spy9                         : std_logic;
  signal srclc                        : std_logic;
  signal srcm                         : std_logic;
  signal srcmap                       : std_logic;
  signal srcmd                        : std_logic;
  signal srcpdlidx                    : std_logic;
  signal srcpdlptr                    : std_logic;
  signal srcq                         : std_logic;
  signal srcvma                       : std_logic;
  signal srun                         : std_logic;
  signal ssdone                       : std_logic;
  signal sspeed0                      : std_logic;
  signal sspeed1                      : std_logic;
  signal sstep                        : std_logic;
  signal st0                          : std_logic;
  signal st10                         : std_logic;
  signal st11                         : std_logic;
  signal st12                         : std_logic;
  signal st13                         : std_logic;
  signal st14                         : std_logic;
  signal st15                         : std_logic;
  signal st16                         : std_logic;
  signal st17                         : std_logic;
  signal st18                         : std_logic;
  signal st19                         : std_logic;
  signal st1                          : std_logic;
  signal st20                         : std_logic;
  signal st21                         : std_logic;
  signal st22                         : std_logic;
  signal st23                         : std_logic;
  signal st24                         : std_logic;
  signal st25                         : std_logic;
  signal st26                         : std_logic;
  signal st27                         : std_logic;
  signal st28                         : std_logic;
  signal st29                         : std_logic;
  signal st2                          : std_logic;
  signal st30                         : std_logic;
  signal st31                         : std_logic;
  signal st3                          : std_logic;
  signal st4                          : std_logic;
  signal st5                          : std_logic;
  signal st6                          : std_logic;
  signal st7                          : std_logic;
  signal st8                          : std_logic;
  signal st9                          : std_logic;
  signal stathenb                     : std_logic;
  signal statstop                     : std_logic;
  signal step                         : std_logic;
  signal tilt0                        : std_logic;
  signal tilt1                        : std_logic;
  signal tpclk                        : std_logic;
  signal tprend                       : std_logic;
  signal tptse                        : std_logic;
  signal tpwp                         : std_logic;
  signal tpwpiram                     : std_logic;
  signal trapa                        : std_logic;
  signal trapb                        : std_logic;
  signal trapenb                      : std_logic;
  signal tse1a                        : std_logic;
  signal tse1b                        : std_logic;
  signal tse2                         : std_logic;
  signal tse3a                        : std_logic;
  signal tse4a                        : std_logic;
  signal tse4b                        : std_logic;
  signal v0parok                      : std_logic;
  signal vcc                          : std_logic;
  signal vm0pari                      : std_logic;
  signal vm1mpar                      : std_logic;
  signal vm1pari                      : std_logic;
  signal vmap0a                       : std_logic;
  signal vmap0b                       : std_logic;
  signal vmap1a                       : std_logic;
  signal vmap1b                       : std_logic;
  signal vmap2a                       : std_logic;
  signal vmap2b                       : std_logic;
  signal vmap3a                       : std_logic;
  signal vmap3b                       : std_logic;
  signal vmap4a                       : std_logic;
  signal vmap4b                       : std_logic;
  signal vmasela                      : std_logic;
  signal vmaselb                      : std_logic;
  signal vmo18                        : std_logic;
  signal vmo19                        : std_logic;
  signal vmopar                       : std_logic;
  signal vmoparck                     : std_logic;
  signal vmoparl                      : std_logic;
  signal vmoparm                      : std_logic;
  signal vmoparodd                    : std_logic;
  signal vmoparok                     : std_logic;
  signal vpari                        : std_logic;
  signal wadr0                        : std_logic;
  signal wadr1                        : std_logic;
  signal wadr2                        : std_logic;
  signal wadr3                        : std_logic;
  signal wadr4                        : std_logic;
  signal wadr5                        : std_logic;
  signal wadr6                        : std_logic;
  signal wadr7                        : std_logic;
  signal wadr8                        : std_logic;
  signal wadr9                        : std_logic;
  signal wmap                         : std_logic;
  signal wmapd                        : std_logic;
  signal wp1a                         : std_logic;
  signal wp1b                         : std_logic;
  signal wp2                          : std_logic;
  signal wp3a                         : std_logic;
  signal wp4a                         : std_logic;
  signal wp4b                         : std_logic;
  signal wp4c                         : std_logic;
  signal wp5a                         : std_logic;
  signal wp5b                         : std_logic;
  signal wp5c                         : std_logic;
  signal wp5d                         : std_logic;
  signal wpc0                         : std_logic;
  signal wpc10                        : std_logic;
  signal wpc11                        : std_logic;
  signal wpc12                        : std_logic;
  signal wpc13                        : std_logic;
  signal wpc1                         : std_logic;
  signal wpc2                         : std_logic;
  signal wpc3                         : std_logic;
  signal wpc4                         : std_logic;
  signal wpc5                         : std_logic;
  signal wpc6                         : std_logic;
  signal wpc7                         : std_logic;
  signal wpc8                         : std_logic;
  signal wpc9                         : std_logic;
  signal wrcyc                        : std_logic;
  signal xout11                       : std_logic;
  signal xout15                       : std_logic;
  signal xout19                       : std_logic;
  signal xout23                       : std_logic;
  signal xout27                       : std_logic;
  signal xout31                       : std_logic;
  signal xout3                        : std_logic;
  signal xout7                        : std_logic;
  signal xx0                          : std_logic;
  signal xx1                          : std_logic;
  signal yout11                       : std_logic;
  signal yout15                       : std_logic;
  signal yout19                       : std_logic;
  signal yout23                       : std_logic;
  signal yout27                       : std_logic;
  signal yout31                       : std_logic;
  signal yout3                        : std_logic;
  signal yout7                        : std_logic;
  signal yy0                          : std_logic;
  signal yy1                          : std_logic;
  signal zero16                       : std_logic;


--- Aliases for some of the above signals to make life easier.

  signal pc : std_logic_vector(0 to 13);  -- Same as PC0, ..., PC13.

begin

  --- Clock Generation

  clock1_1c08 : ic_74s10 port map(g1a   => \-clock_reset_b\, g1b => \-tpdone\, g2a=>\-hang\, g2b=>\-clock_reset_b\, g2c=>cyclecompleted, g2y_n=>\-tpr0\, g1y_n=>internal12, g1c=>internal11, g3a=>'0', g3b=>'0', g3c=>'0');
  clock1_1c09 : ic_74s00 port map(g1b   => internal12, g1a => \-tpr40\, g1q_n => internal11, g2b => '0', g2a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  clock1_1c10 : ic_74s02 port map(g4b   => internal11, g4a => gnd, g4q_n => cyclecompleted, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g3b => '0', g3a => '0');
  clock1_1c12 : ic_td50 port map(input  => \-tprend\, o_20ns => \-tpw20\, o_40ns=>\-tpw40\, o_50ns=>\-tpw50\, o_30ns=>\-tpw30\, o_10ns=>\-tpw10\);
  clock1_1c14 : ic_td25 port map(input  => \-tpw50\, o_10ns => \-tpw60\, o_20ns=>\-tpw70\, o_25ns=>\-tpw75\, o_15ns=>\-tpw65\, o_5ns=>\-tpw55\);
  clock1_1c15 : ic_td25 port map(input  => \-tpw20\, o_10ns => \-tpw30a\, o_20ns=>\-tpw40a\, o_25ns=>\-tpw45\, o_15ns=>\-tpw35\, o_5ns=>\-tpw25\);
  clock1_1d08 : ic_74s151 port map(i3   => \-tpr100\, i2 => \-tpr140\, i1=>\-tpr160\, i0=>\-tpr160\, q=>\-tprend\, q_n=>tprend, ce_n=>gnd, sel2=>sspeed1, sel1=>sspeed0, sel0=>\-ilong\, i7=>\-tpr75\, i6=>\-tpr115\, i5=>\-tpr85\, i4=>\-tpr125\);
  clock1_1d11 : ic_td25 port map(input  => \-tpr0\, o_10ns => \-tpr10\, o_20ns=>\-tpr20a\, o_25ns=>\-tpr25\, o_15ns=>\-tpr15\, o_5ns=>\-tpr5\);
  clock1_1d12 : ic_td100 port map(input => \-tpr0\, o_40ns => \-tpr40\, o_80ns=>\-tpr80\, o_100ns=>\-tpr100\, o_60ns=>\-tpr60\, o_20ns=>\-tpr20\);
  clock1_1d13 : ic_td100 port map(input => \-tpr100\, o_40ns => \-tpr140\, o_80ns=>\-tpr180\, o_100ns=>\-tpr200\, o_60ns=>\-tpr160\, o_20ns=>\-tpr120\);
  clock1_1d14 : ic_td25 port map(input  => \-tpr100\, o_10ns => \-tpr110\, o_20ns=>\-tpr120a\, o_25ns=>\-tpr125\, o_15ns=>\-tpr115\, o_5ns=>\-tpr105\);
  clock1_1d15 : ic_td25 port map(input  => \-tpr60\, o_10ns => \-tpr70\, o_20ns=>\-tpr80a\, o_25ns=>\-tpr85\, o_15ns=>\-tpr75\, o_5ns=>\-tpr65\);

  clock2_1c01 : ic_7428 port map(g1q_n  => clk4, g1a => \-clk0\, g1b => gnd, g2q_n => mclk7, g2a => \-mclk0\, g2b=>gnd, g3a=>'0', g4a=>'0', g4b=>'0', g3b=>'0');
  clock2_1c02 : ic_7428 port map(g1q_n  => \-wp1\, g1a => tpwp, g1b => gnd, g2q_n => \-wp2\, g2a=>tpwp, g2b=>gnd, g3a=>gnd, g3b=>tpwp, g3q_n=>\-wp3\, g4a=>gnd, g4b=>tpwp, g4q_n=>\-wp4\);
  clock2_1c06 : ic_74s10 port map(g1a   => \-tprend\, g1b => tpclk, g2a => \-tptse\, g2b=>\-tpr25\, g2c=>\-clock_reset_b\, g2y_n=>tptse, g3y_n=>internal7, g3a=>\-clock_reset_b\, g3b=>\-tpw70\, g3c=>internal10, g1y_n=>\-tpclk\, g1c=>\-clock_reset_b\);
  clock2_1c07 : ic_74s00 port map(g1b   => \-tpr0\, g1a => \-tpclk\, g1q_n=>tpclk, g2b=>\-tpr5\, g2a=>tptse, g2q_n=>\-tptse\, g3q_n=>internal10, g3b=>internal7, g3a=>\-tpw30\, g4a=>'0', g4b=>'0');
  clock2_1c10 : ic_74s02 port map(g2q_n => tpwp, g2a => internal7, g2b => \machruna_l\, g3b => \machruna_l\, g3a=>internal8, g3q_n=>tpwpiram, g1a=>'0', g1b=>'0', g4b=>'0', g4a=>'0');
  clock2_1c11 : ic_7428 port map(g1q_n  => \-wp5\, g1a => tpwpiram, g1b => gnd, g2q_n => clk5, g2a => \-clk0\, g2b=>gnd, g3a=>gnd, g3b=>\-mclk0\, g3q_n=>mclk5, g4a=>'0', g4b=>'0');
  clock2_1c13 : ic_74s10 port map(g2a   => \-tprend\, g2b => internal8, g2c => internal8, g2y_n => internal9, g3y_n => internal8, g3a => \-tpw45\, g3b=>\-clock_reset_b\, g3c=>internal9, g1a=>'0', g1b=>'0', g1c=>'0');
  clock2_1d04 : ic_7428 port map(g1q_n  => \-tse1\, g1a => tptse, g1b => gnd, g2q_n => \-tse2\, g2a=>tptse, g2b=>gnd, g3a=>gnd, g3b=>tptse, g3q_n=>\-tse3\, g4a=>gnd, g4b=>tptse, g4q_n=>\-tse4\);
  clock2_1d05 : ic_7428 port map(g1q_n  => clk1, g1a => \-clk0\, g1b => gnd, g2q_n => clk2, g2a => \-clk0\, g2b=>gnd, g3a=>gnd, g3b=>\-clk0\, g3q_n=>clk3, g4a=>gnd, g4b=>\-mclk0\, g4q_n=>mclk1);
  clock2_1d10 : ic_74s08 port map(g1b   => \-tpclk\, g1a => machrun, g1q => \-clk0\, g3q=>\-mclk0\, g3a=>hi1, g3b=>\-tpclk\, g2b=>'0', g2a=>'0', g4a=>'0', g4b=>'0');

  clockd_1b18 : ic_74s37 port map(g1a => \-clk1\, g1b => hi12, g1y => clk1a, g2a => reset, g2b => hi12, g2y => \-reset\, g3y=>mclk1a, g3a=>hi12, g3b=>\-mclk1\, g4a=>'0', g4b=>'0');
  clockd_1b19 : ic_74s04 port map(g1a => mclk1, g1q_n => \-mclk1\, g2a => clk1, g2q_n => \-clk1\, g3a=>\-wp1\, g3q_n=>wp1b, g4q=>wp1a, g4a=>\-wp1\, g5q_n=>tse1b, g5a=>\-tse1\, g6q_n=>tse1a, g6a=>\-tse1\);
  clockd_1f05 : ic_74s133 port map(g  => hi1, f => hi2, e => hi3, d => hi4, c => hi5, b => hi6, a => hi7, q_n => \-upperhighok\, h => hi8, i => hi9, j => hi10, k => hi11, l => hi12, m => hi11);
  clockd_2c02 : ic_74s04 port map(g1a => lcry3, g1q_n => \-lcry3\, g2a => nc429, g2q_n => nc430, g3a => clk2, g3q_n => \-clk2c\, g4q=>\-clk2a\, g4a=>clk2, g5q_n=>wp2, g5a=>\-wp2\, g6q_n=>tse2, g6a=>\-tse2\);
  clockd_2c03 : ic_74s37 port map(g1a => \-clk2a\, g1b => hi7, g1y => clk2a, g2a => \-clk2a\, g2b=>hi7, g2y=>clk2b, g3y=>clk2c, g3a=>hi7, g3b=>\-clk2c\, g4a=>'0', g4b=>'0');
  clockd_3c11 : ic_74s37 port map(g1a => \-clk3a\, g1b => hi5, g1y => clk3a, g2a => \-clk3a\, g2b=>hi5, g2y=>clk3b, g3y=>clk3c, g3a=>hi5, g3b=>\-clk3a\, g4a=>'0', g4b=>'0');
  clockd_3c12 : ic_74s04 port map(g1a => nc427, g1q_n => nc428, g2a => clk3, g2q_n => \-clk3g\, g3a => clk3, g3q_n => \-clk3d\, g4q=>\-clk3a\, g4a=>clk3, g5q_n=>wp3a, g5a=>\-wp3\, g6q_n=>tse3a, g6a=>\-tse3\);
  clockd_3c13 : ic_74s37 port map(g1a => \-clk3d\, g1b => hi5, g1y => clk3d, g2a => \-clk3d\, g2b=>hi5, g2y=>clk3e, g3y=>clk3f, g3a=>hi5, g3b=>\-clk3d\, g4a=>'0', g4b=>'0');
  clockd_4c02 : ic_74s37 port map(g1a => \-clk4a\, g1b => hi5, g1y => clk4a, g2a => \-clk4a\, g2b=>hi5, g2y=>clk4b, g3y=>clk4c, g3a=>hi5, g3b=>\-clk4a\, g4a=>'0', g4b=>'0');
  clockd_4c06 : ic_74s04 port map(g1a => clk4, g1q_n => \-clk4e\, g2a => clk4, g2q_n => \-clk4d\, g3a=>clk4, g3q_n=>\-clk4a\, g4q=>wp4c, g4a=>\-wp4\, g5q_n=>wp4b, g5a=>\-wp4\, g6q_n=>wp4a, g6a=>\-wp4\);
  clockd_4c07 : ic_74s37 port map(g1a => \-clk4d\, g1b => hi2, g1y => clk4d, g2a => \-clk4d\, g2b=>hi2, g2y=>clk4e, g3y=>clk4f, g3a=>hi2, g3b=>\-clk4d\, g4a=>'0', g4b=>'0');
  clockd_4d03 : ic_74s04 port map(g1a => nc423, g1q_n => nc424, g2a => nc425, g2q_n => nc426, g3a => \-tse4\, g3q_n => tse4b, g4q => tse4a, g4a => \-tse4\, g5q_n=>srcpdlptr, g5a=>\-srcpdlptr\, g6q_n=>srcpdlidx, g6a=>\-srcpdlidx\);

  --- Microinstruction Fetch

  ictl_1a15 : ic_9s42_1 port map(out2 => ramdisable, g2d2 => hi1, g2c2 => hi1, g2b2 => \-iwriteda\, g2a2 => \-promdisabled\, g1b2=>hi1, g1a2=>idebug, g1a1=>'0', g1b1=>'0', g2a1=>'0', g2b1=>'0', g2c1=>'0', g2d1=>'0');
  ictl_1c16 : ic_74s04 port map(g1a   => iwriteda, g1q_n => \-iwriteda\, g2a => promdisabled, g2q_n => \-promdisabled\, g3a=>\-wp5\, g3q_n=>wp5d, g4q=>wp5c, g4a=>\-wp5\, g5q_n=>wp5b, g5a=>\-wp5\, g6q_n=>wp5a, g6a=>\-wp5\);
  ictl_1c21 : ic_74s04 port map(g1a   => pc0, g1q_n => \-pcb0\, g2a => pc1, g2q_n => \-pcb1\, g3a=>pc2, g3q_n=>\-pcb2\, g4q=>\-pcb3\, g4a=>pc3, g5q_n=>\-pcb4\, g5a=>pc4, g6q_n=>\-pcb5\, g6a=>pc5);
  ictl_1c26 : ic_74s37 port map(g1a   => wp5a, g1b => iwriteda, g1y => \-iwea\, g2a => wp5a, g2b => iwriteda, g2y => \-iweb\, g3y=>\-iwei\, g3a=>iwriteda, g3b=>wp5a, g4y=>\-iwej\, g4a=>iwriteda, g4b=>wp5a);
  ictl_1d20 : ic_74s04 port map(g1a   => pc13, g1q_n => \-pc13b\, g2a => pc12, g2q_n => \-pc12b\, g3a=>\-iwrited\, g3q_n=>iwritedd, g4q=>iwritedc, g4a=>\-iwrited\, g5q_n=>iwritedb, g5a=>\-iwrited\, g6q_n=>iwriteda, g6a=>\-iwrited\);
  ictl_1d25 : ic_74s04 port map(g1a   => pc6, g1q_n => \-pcb6\, g2a => pc7, g2q_n => \-pcb7\, g3a=>pc8, g3q_n=>\-pcb8\, g4q=>\-pcb9\, g4a=>pc9, g5q_n=>\-pcb10\, g5a=>pc10, g6q_n=>\-pcb11\, g6a=>pc11);
  ictl_1d30 : ic_74s139 port map(g1   => ramdisable, a1 => \-pc12b\, b1 => \-pc13b\, g1y0=>\-ice3a\, g1y1=>\-ice2a\, g1y2=>\-ice1a\, g1y3=>\-ice0a\, g2y3=>\-ice0b\, g2y2=>\-ice1b\, g2y1=>\-ice2b\, g2y0=>\-ice3b\, b2=>\-pc13b\, a2=>\-pc12b\, g2=>ramdisable);
  ictl_2c01 : ic_74s37 port map(g1a   => wp5b, g1b => iwritedb, g1y => \-iwec\, g2a => wp5b, g2b => iwritedb, g2y => \-iwed\, g3y=>\-iwek\, g3a=>iwritedb, g3b=>wp5b, g4y=>\-iwel\, g4a=>iwritedb, g4b=>wp5b);
  ictl_2c06 : ic_74s04 port map(g1a   => pc0, g1q_n => \-pcc0\, g2a => pc1, g2q_n => \-pcc1\, g3a=>pc2, g3q_n=>\-pcc2\, g4q=>\-pcc3\, g4a=>pc3, g5q_n=>\-pcc4\, g5a=>pc4, g6q_n=>\-pcc5\, g6a=>pc5);
  ictl_2d10 : ic_74s04 port map(g1a   => pc6, g1q_n => \-pcc6\, g2a => pc7, g2q_n => \-pcc7\, g3a=>pc8, g3q_n=>\-pcc8\, g4q=>\-pcc9\, g4a=>pc9, g5q_n=>\-pcc10\, g5a=>pc10, g6q_n=>\-pcc11\, g6a=>pc11);
  ictl_2d15 : ic_74s37 port map(g1a   => wp5c, g1b => iwritedc, g1y => \-iwee\, g2a => wp5c, g2b => iwritedc, g2y => \-iwef\, g3y=>\-iwem\, g3a=>iwritedc, g3b=>wp5c, g4y=>\-iwen\, g4a=>iwritedc, g4b=>wp5c);
  ictl_2d25 : ic_74s139 port map(g1   => ramdisable, a1 => \-pc12b\, b1 => \-pc13b\, g1y0=>\-ice3c\, g1y1=>\-ice2c\, g1y2=>\-ice1c\, g1y3=>\-ice0c\, g2y3=>\-ice0d\, g2y2=>\-ice1d\, g2y1=>\-ice2d\, g2y0=>\-ice3d\, b2=>\-pc13b\, a2=>\-pc12b\, g2=>ramdisable);
  ictl_2d30 : ic_74s37 port map(g1a   => wp5d, g1b => iwritedd, g1y => \-iweg\, g2a => wp5d, g2b => iwritedd, g2y => \-iweh\, g3y=>\-iweo\, g3a=>iwritedd, g3b=>wp5d, g4y=>\-iwep\, g4a=>iwritedd, g4b=>wp5d);

  iram00_1d21 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i10, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr10, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1d22 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i11, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr11, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1d23 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6a, g2a => \-pcb7\, g2q_n=>pc7a, g3a=>\-pcb8\, g3q_n=>pc8a, g4q=>pc9a, g4a=>\-pcb9\, g5q_n=>pc10a, g5a=>\-pcb10\, g6q_n=>pc11a, g6a=>\-pcb11\);
  iram00_1d24 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0a, g2a => \-pcb1\, g2q_n=>pc1a, g3a=>\-pcb2\, g3q_n=>pc2a, g4q=>pc3a, g4a=>\-pcb3\, g5q_n=>pc4a, g5a=>\-pcb4\, g6q_n=>pc5a, g6a=>\-pcb5\);
  iram00_1e21 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i5, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr5, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1e22 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i6, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr6, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1e23 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i7, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr7, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1e24 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i8, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr8, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1e25 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i9, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr9, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1f21 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i0, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr0, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1f22 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i1, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr1, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1f23 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i2, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr2, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1f24 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i3, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr3, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);
  iram00_1f25 : ic_2147 port map(a0   => pc0a, a1 => pc1a, a2 => pc2a, a3 => pc3a, a4 => pc4a, a5 => pc5a, do => i4, we_n => \-iwea\, ce_n => \-ice0a\, di=>iwr4, a11=>pc11a, a10=>pc10a, a9=>pc9a, a8=>pc8a, a7=>pc7a, a6=>pc6a);

  iram01_1d26 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i10, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr10, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1d27 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i11, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr11, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1d28 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6b, g2a => \-pcb7\, g2q_n=>pc7b, g3a=>\-pcb8\, g3q_n=>pc8b, g4q=>pc9b, g4a=>\-pcb9\, g5q_n=>pc10b, g5a=>\-pcb10\, g6q_n=>pc11b, g6a=>\-pcb11\);
  iram01_1d29 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0b, g2a => \-pcb1\, g2q_n=>pc1b, g3a=>\-pcb2\, g3q_n=>pc2b, g4q=>pc3b, g4a=>\-pcb3\, g5q_n=>pc4b, g5a=>\-pcb4\, g6q_n=>pc5b, g6a=>\-pcb5\);
  iram01_1e26 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i5, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr5, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1e27 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i6, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr6, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1e28 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i7, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr7, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1e29 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i8, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr8, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1e30 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i9, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr9, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1f26 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i0, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr0, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1f27 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i1, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr1, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1f28 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i2, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr2, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1f29 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i3, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr3, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);
  iram01_1f30 : ic_2147 port map(a0   => pc0b, a1 => pc1b, a2 => pc2b, a3 => pc3b, a4 => pc4b, a5 => pc5b, do => i4, we_n => \-iweb\, ce_n => \-ice1a\, di=>iwr4, a11=>pc11b, a10=>pc10b, a9=>pc9b, a8=>pc8b, a7=>pc7b, a6=>pc6b);

  iram02_2d01 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i10, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr10, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2d02 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i11, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr11, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2d03 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6c, g2a => \-pcb7\, g2q_n=>pc7c, g3a=>\-pcb8\, g3q_n=>pc8c, g4q=>pc9c, g4a=>\-pcb9\, g5q_n=>pc10c, g5a=>\-pcb10\, g6q_n=>pc11c, g6a=>\-pcb11\);
  iram02_2d04 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0c, g2a => \-pcb1\, g2q_n=>pc1c, g3a=>\-pcb2\, g3q_n=>pc2c, g4q=>pc3c, g4a=>\-pcb3\, g5q_n=>pc4c, g5a=>\-pcb4\, g6q_n=>pc5c, g6a=>\-pcb5\);
  iram02_2e01 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i5, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr5, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2e02 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i6, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr6, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2e03 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i7, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr7, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2e04 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i8, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr8, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2e05 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i9, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr9, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2f01 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i0, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr0, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2f02 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i1, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr1, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2f03 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i2, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr2, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2f04 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i3, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr3, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);
  iram02_2f05 : ic_2147 port map(a0   => pc0c, a1 => pc1c, a2 => pc2c, a3 => pc3c, a4 => pc4c, a5 => pc5c, do => i4, we_n => \-iwec\, ce_n => \-ice2a\, di=>iwr4, a11=>pc11c, a10=>pc10c, a9=>pc9c, a8=>pc8c, a7=>pc7c, a6=>pc6c);

  iram03_2d06 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i10, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr10, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2d07 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i11, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr11, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2d08 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6d, g2a => \-pcb7\, g2q_n=>pc7d, g3a=>\-pcb8\, g3q_n=>pc8d, g4q=>pc9d, g4a=>\-pcb9\, g5q_n=>pc10d, g5a=>\-pcb10\, g6q_n=>pc11d, g6a=>\-pcb11\);
  iram03_2d09 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0d, g2a => \-pcb1\, g2q_n=>pc1d, g3a=>\-pcb2\, g3q_n=>pc2d, g4q=>pc3d, g4a=>\-pcb3\, g5q_n=>pc4d, g5a=>\-pcb4\, g6q_n=>pc5d, g6a=>\-pcb5\);
  iram03_2e06 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i5, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr5, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2e07 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i6, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr6, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2e08 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i7, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr7, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2e09 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i8, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr8, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2e10 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i9, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr9, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2f06 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i0, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr0, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2f07 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i1, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr1, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2f08 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i2, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr2, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2f09 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i3, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr3, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);
  iram03_2f10 : ic_2147 port map(a0   => pc0d, a1 => pc1d, a2 => pc2d, a3 => pc3d, a4 => pc4d, a5 => pc5d, do => i4, we_n => \-iwed\, ce_n => \-ice3a\, di=>iwr4, a11=>pc11d, a10=>pc10d, a9=>pc9d, a8=>pc8d, a7=>pc7d, a6=>pc6d);

  iram10_2d11 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i22, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr22, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2d12 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i23, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr23, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2d13 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6e, g2a => \-pcb7\, g2q_n=>pc7e, g3a=>\-pcb8\, g3q_n=>pc8e, g4q=>pc9e, g4a=>\-pcb9\, g5q_n=>pc10e, g5a=>\-pcb10\, g6q_n=>pc11e, g6a=>\-pcb11\);
  iram10_2d14 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0e, g2a => \-pcb1\, g2q_n=>pc1e, g3a=>\-pcb2\, g3q_n=>pc2e, g4q=>pc3e, g4a=>\-pcb3\, g5q_n=>pc4e, g5a=>\-pcb4\, g6q_n=>pc5e, g6a=>\-pcb5\);
  iram10_2e11 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i17, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr17, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2e12 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i18, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr18, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2e13 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i19, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr19, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2e14 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i20, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr20, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2e15 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i21, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr21, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2f11 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i12, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr12, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2f12 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i13, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr13, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2f13 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i14, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr14, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2f14 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i15, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr15, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);
  iram10_2f15 : ic_2147 port map(a0   => pc0e, a1 => pc1e, a2 => pc2e, a3 => pc3e, a4 => pc4e, a5 => pc5e, do => i16, we_n => \-iwee\, ce_n => \-ice0b\, di=>iwr16, a11=>pc11e, a10=>pc10e, a9=>pc9e, a8=>pc8e, a7=>pc7e, a6=>pc6e);

  iram11_2d16 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i22, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr22, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2d17 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i23, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr23, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2d18 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6f, g2a => \-pcb7\, g2q_n=>pc7f, g3a=>\-pcb8\, g3q_n=>pc8f, g4q=>pc9f, g4a=>\-pcb9\, g5q_n=>pc10f, g5a=>\-pcb10\, g6q_n=>pc11f, g6a=>\-pcb11\);
  iram11_2d19 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0f, g2a => \-pcb1\, g2q_n=>pc1f, g3a=>\-pcb2\, g3q_n=>pc2f, g4q=>pc3f, g4a=>\-pcb3\, g5q_n=>pc4f, g5a=>\-pcb4\, g6q_n=>pc5f, g6a=>\-pcb5\);
  iram11_2e16 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i17, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr17, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2e17 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i18, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr18, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2e18 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i19, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr19, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2e19 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i20, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr20, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2e20 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i21, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr21, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2f16 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i12, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr12, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2f17 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i13, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr13, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2f18 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i14, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr14, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2f19 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i15, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr15, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);
  iram11_2f20 : ic_2147 port map(a0   => pc0f, a1 => pc1f, a2 => pc2f, a3 => pc3f, a4 => pc4f, a5 => pc5f, do => i16, we_n => \-iwef\, ce_n => \-ice1b\, di=>iwr16, a11=>pc11f, a10=>pc10f, a9=>pc9f, a8=>pc8f, a7=>pc7f, a6=>pc6f);

  iram12_2d21 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i22, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr22, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2d22 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i23, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr23, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2d23 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6g, g2a => \-pcb7\, g2q_n=>pc7g, g3a=>\-pcb8\, g3q_n=>pc8g, g4q=>pc9g, g4a=>\-pcb9\, g5q_n=>pc10g, g5a=>\-pcb10\, g6q_n=>pc11g, g6a=>\-pcb11\);
  iram12_2d24 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0g, g2a => \-pcb1\, g2q_n=>pc1g, g3a=>\-pcb2\, g3q_n=>pc2g, g4q=>pc3g, g4a=>\-pcb3\, g5q_n=>pc4g, g5a=>\-pcb4\, g6q_n=>pc5g, g6a=>\-pcb5\);
  iram12_2e21 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i17, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr17, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2e22 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i18, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr18, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2e23 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i19, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr19, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2e24 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i20, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr20, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2e25 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i21, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr21, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2f21 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i12, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr12, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2f22 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i13, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr13, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2f23 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i14, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr14, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2f24 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i15, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr15, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);
  iram12_2f25 : ic_2147 port map(a0   => pc0g, a1 => pc1g, a2 => pc2g, a3 => pc3g, a4 => pc4g, a5 => pc5g, do => i16, we_n => \-iweg\, ce_n => \-ice2b\, di=>iwr16, a11=>pc11g, a10=>pc10g, a9=>pc9g, a8=>pc8g, a7=>pc7g, a6=>pc6g);

  iram13_2d26 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i22, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr22, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2d27 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i23, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr23, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2d28 : ic_74s04 port map(g1a => \-pcb6\, g1q_n => pc6h, g2a => \-pcb7\, g2q_n=>pc7h, g3a=>\-pcb8\, g3q_n=>pc8h, g4q=>pc9h, g4a=>\-pcb9\, g5q_n=>pc10h, g5a=>\-pcb10\, g6q_n=>pc11h, g6a=>\-pcb11\);
  iram13_2d29 : ic_74s04 port map(g1a => \-pcb0\, g1q_n => pc0h, g2a => \-pcb1\, g2q_n=>pc1h, g3a=>\-pcb2\, g3q_n=>pc2h, g4q=>pc3h, g4a=>\-pcb3\, g5q_n=>pc4h, g5a=>\-pcb4\, g6q_n=>pc5h, g6a=>\-pcb5\);
  iram13_2e26 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i17, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr17, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2e27 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i18, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr18, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2e28 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i19, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr19, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2e29 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i20, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr20, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2e30 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i21, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr21, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2f26 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i12, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr12, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2f27 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i13, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr13, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2f28 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i14, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr14, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2f29 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i15, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr15, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);
  iram13_2f30 : ic_2147 port map(a0   => pc0h, a1 => pc1h, a2 => pc2h, a3 => pc3h, a4 => pc4h, a5 => pc5h, do => i16, we_n => \-iweh\, ce_n => \-ice3b\, di=>iwr16, a11=>pc11h, a10=>pc10h, a9=>pc9h, a8=>pc8h, a7=>pc7h, a6=>pc6h);

  iram20_1a21 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i31, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr31, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1a22 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i32, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr32, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1a23 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i33, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr33, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1a24 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i34, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr34, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1a25 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i35, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr35, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1b21 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i26, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr26, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1b22 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i27, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr27, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1b23 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i28, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr28, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1b24 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i29, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr29, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1b25 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i30, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr30, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1c22 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6i, g2a => \-pcc7\, g2q_n=>pc7i, g3a=>\-pcc8\, g3q_n=>pc8i, g4q=>pc9i, g4a=>\-pcc9\, g5q_n=>pc10i, g5a=>\-pcc10\, g6q_n=>pc11i, g6a=>\-pcc11\);
  iram20_1c23 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0i, g2a => \-pcc1\, g2q_n=>pc1i, g3a=>\-pcc2\, g3q_n=>pc2i, g4q=>pc3i, g4a=>\-pcc3\, g5q_n=>pc4i, g5a=>\-pcc4\, g6q_n=>pc5i, g6a=>\-pcc5\);
  iram20_1c24 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i24, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr24, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);
  iram20_1c25 : ic_2147 port map(a0   => pc0i, a1 => pc1i, a2 => pc2i, a3 => pc3i, a4 => pc4i, a5 => pc5i, do => i25, we_n => \-iwei\, ce_n => \-ice0c\, di=>iwr25, a11=>pc11i, a10=>pc10i, a9=>pc9i, a8=>pc8i, a7=>pc7i, a6=>pc6i);

  iram21_1a26 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i31, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr31, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1a27 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i32, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr32, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1a28 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i33, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr33, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1a29 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i34, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr34, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1a30 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i35, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr35, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1b26 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i26, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr26, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1b27 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i27, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr27, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1b28 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i28, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr28, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1b29 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i29, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr29, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1b30 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i30, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr30, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1c27 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6j, g2a => \-pcc7\, g2q_n=>pc7j, g3a=>\-pcc8\, g3q_n=>pc8j, g4q=>pc9j, g4a=>\-pcc9\, g5q_n=>pc10j, g5a=>\-pcc10\, g6q_n=>pc11j, g6a=>\-pcc11\);
  iram21_1c28 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0j, g2a => \-pcc1\, g2q_n=>pc1j, g3a=>\-pcc2\, g3q_n=>pc2j, g4q=>pc3j, g4a=>\-pcc3\, g5q_n=>pc4j, g5a=>\-pcc4\, g6q_n=>pc5j, g6a=>\-pcc5\);
  iram21_1c29 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i24, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr24, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);
  iram21_1c30 : ic_2147 port map(a0   => pc0j, a1 => pc1j, a2 => pc2j, a3 => pc3j, a4 => pc4j, a5 => pc5j, do => i25, we_n => \-iwej\, ce_n => \-ice1c\, di=>iwr25, a11=>pc11j, a10=>pc10j, a9=>pc9j, a8=>pc8j, a7=>pc7j, a6=>pc6j);

  iram22_2a01 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i31, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr31, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2a02 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i32, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr32, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2a03 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i33, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr33, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2a04 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i34, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr34, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2a05 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i35, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr35, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2b01 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i26, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr26, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2b02 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i27, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr27, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2b03 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i28, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr28, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2b04 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i29, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr29, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2b05 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i30, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr30, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2c02 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6k, g2a => \-pcc7\, g2q_n=>pc7k, g3a=>\-pcc8\, g3q_n=>pc8k, g4q=>pc9k, g4a=>\-pcc9\, g5q_n=>pc10k, g5a=>\-pcc10\, g6q_n=>pc11k, g6a=>\-pcc11\);
  iram22_2c03 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0k, g2a => \-pcc1\, g2q_n=>pc1k, g3a=>\-pcc2\, g3q_n=>pc2k, g4q=>pc3k, g4a=>\-pcc3\, g5q_n=>pc4k, g5a=>\-pcc4\, g6q_n=>pc5k, g6a=>\-pcc5\);
  iram22_2c04 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i24, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr24, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);
  iram22_2c05 : ic_2147 port map(a0   => pc0k, a1 => pc1k, a2 => pc2k, a3 => pc3k, a4 => pc4k, a5 => pc5k, do => i25, we_n => \-iwek\, ce_n => \-ice2c\, di=>iwr25, a11=>pc11k, a10=>pc10k, a9=>pc9k, a8=>pc8k, a7=>pc7k, a6=>pc6k);

  iram23_2a06 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i31, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr31, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2a07 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i32, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr32, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2a08 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i33, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr33, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2a09 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i34, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr34, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2a10 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i35, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr35, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2b06 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i26, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr26, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2b07 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i27, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr27, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2b08 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i28, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr28, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2b09 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i29, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr29, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2b10 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i30, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr30, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2c07 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6l, g2a => \-pcc7\, g2q_n=>pc7l, g3a=>\-pcc8\, g3q_n=>pc8l, g4q=>pc9l, g4a=>\-pcc9\, g5q_n=>pc10l, g5a=>\-pcc10\, g6q_n=>pc11l, g6a=>\-pcc11\);
  iram23_2c08 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0l, g2a => \-pcc1\, g2q_n=>pc1l, g3a=>\-pcc2\, g3q_n=>pc2l, g4q=>pc3l, g4a=>\-pcc3\, g5q_n=>pc4l, g5a=>\-pcc4\, g6q_n=>pc5l, g6a=>\-pcc5\);
  iram23_2c09 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i24, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr24, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);
  iram23_2c10 : ic_2147 port map(a0   => pc0l, a1 => pc1l, a2 => pc2l, a3 => pc3l, a4 => pc4l, a5 => pc5l, do => i25, we_n => \-iwel\, ce_n => \-ice3c\, di=>iwr25, a11=>pc11l, a10=>pc10l, a9=>pc9l, a8=>pc8l, a7=>pc7l, a6=>pc6l);

  iram30_2a11 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i44, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr44, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2a12 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i45, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr45, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2a13 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i46, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr46, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2a14 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i47, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr47, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2a15 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i48, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr48, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2b11 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i39, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr39, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2b12 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i40, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr40, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2b13 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i41, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr41, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2b14 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i42, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr42, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2b15 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i43, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr43, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2c11 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6m, g2a => \-pcc7\, g2q_n=>pc7m, g3a=>\-pcc8\, g3q_n=>pc8m, g4q=>pc9m, g4a=>\-pcc9\, g5q_n=>pc10m, g5a=>\-pcc10\, g6q_n=>pc11m, g6a=>\-pcc11\);
  iram30_2c12 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0m, g2a => \-pcc1\, g2q_n=>pc1m, g3a=>\-pcc2\, g3q_n=>pc2m, g4q=>pc3m, g4a=>\-pcc3\, g5q_n=>pc4m, g5a=>\-pcc4\, g6q_n=>pc5m, g6a=>\-pcc5\);
  iram30_2c13 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i36, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr36, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2c14 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i37, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr37, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);
  iram30_2c15 : ic_2147 port map(a0   => pc0m, a1 => pc1m, a2 => pc2m, a3 => pc3m, a4 => pc4m, a5 => pc5m, do => i38, we_n => \-iwem\, ce_n => \-ice0d\, di=>iwr38, a11=>pc11m, a10=>pc10m, a9=>pc9m, a8=>pc8m, a7=>pc7m, a6=>pc6m);

  iram31_2a16 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i44, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr44, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2a17 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i45, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr45, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2a18 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i46, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr46, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2a19 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i47, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr47, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2a20 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i48, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr48, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2b16 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i39, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr39, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2b17 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i40, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr40, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2b18 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i41, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr41, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2b19 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i42, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr42, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2b20 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i43, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr43, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2c16 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6n, g2a => \-pcc7\, g2q_n=>pc7n, g3a=>\-pcc8\, g3q_n=>pc8n, g4q=>pc9n, g4a=>\-pcc9\, g5q_n=>pc10n, g5a=>\-pcc10\, g6q_n=>pc11n, g6a=>\-pcc11\);
  iram31_2c17 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0n, g2a => \-pcc1\, g2q_n=>pc1n, g3a=>\-pcc2\, g3q_n=>pc2n, g4q=>pc3n, g4a=>\-pcc3\, g5q_n=>pc4n, g5a=>\-pcc4\, g6q_n=>pc5n, g6a=>\-pcc5\);
  iram31_2c18 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i36, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr36, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2c19 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i37, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr37, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);
  iram31_2c20 : ic_2147 port map(a0   => pc0n, a1 => pc1n, a2 => pc2n, a3 => pc3n, a4 => pc4n, a5 => pc5n, do => i38, we_n => \-iwen\, ce_n => \-ice1d\, di=>iwr38, a11=>pc11n, a10=>pc10n, a9=>pc9n, a8=>pc8n, a7=>pc7n, a6=>pc6n);

  iram32_2a21 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i44, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr44, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2a22 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i45, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr45, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2a23 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i46, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr46, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2a24 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i47, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr47, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2a25 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i48, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr48, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2b21 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i39, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr39, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2b22 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i40, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr40, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2b23 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i41, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr41, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2b24 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i42, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr42, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2b25 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i43, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr43, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2c21 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6o, g2a => \-pcc7\, g2q_n=>pc7o, g3a=>\-pcc8\, g3q_n=>pc8o, g4q=>pc9o, g4a=>\-pcc9\, g5q_n=>pc10o, g5a=>\-pcc10\, g6q_n=>pc11o, g6a=>\-pcc11\);
  iram32_2c22 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0o, g2a => \-pcc1\, g2q_n=>pc1o, g3a=>\-pcc2\, g3q_n=>pc2o, g4q=>pc3o, g4a=>\-pcc3\, g5q_n=>pc4o, g5a=>\-pcc4\, g6q_n=>pc5o, g6a=>\-pcc5\);
  iram32_2c23 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i36, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr36, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2c24 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i37, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr37, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);
  iram32_2c25 : ic_2147 port map(a0   => pc0o, a1 => pc1o, a2 => pc2o, a3 => pc3o, a4 => pc4o, a5 => pc5o, do => i38, we_n => \-iweo\, ce_n => \-ice2d\, di=>iwr38, a11=>pc11o, a10=>pc10o, a9=>pc9o, a8=>pc8o, a7=>pc7o, a6=>pc6o);

  iram33_2a26 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i44, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr44, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2a27 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i45, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr45, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2a28 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i46, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr46, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2a29 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i47, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr47, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2a30 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i48, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr48, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2b26 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i39, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr39, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2b27 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i40, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr40, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2b28 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i41, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr41, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2b29 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i42, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr42, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2b30 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i43, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr43, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2c26 : ic_74s04 port map(g1a => \-pcc6\, g1q_n => pc6p, g2a => \-pcc7\, g2q_n=>pc7p, g3a=>\-pcc8\, g3q_n=>pc8p, g4q=>pc9p, g4a=>\-pcc9\, g5q_n=>pc10p, g5a=>\-pcc10\, g6q_n=>pc11p, g6a=>\-pcc11\);
  iram33_2c27 : ic_74s04 port map(g1a => \-pcc0\, g1q_n => pc0p, g2a => \-pcc1\, g2q_n=>pc1p, g3a=>\-pcc2\, g3q_n=>pc2p, g4q=>pc3p, g4a=>\-pcc3\, g5q_n=>pc4p, g5a=>\-pcc4\, g6q_n=>pc5p, g6a=>\-pcc5\);
  iram33_2c28 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i36, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr36, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2c29 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i37, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr37, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);
  iram33_2c30 : ic_2147 port map(a0   => pc0p, a1 => pc1p, a2 => pc2p, a3 => pc3p, a4 => pc4p, a5 => pc5p, do => i38, we_n => \-iwep\, ce_n => \-ice3d\, di=>iwr38, a11=>pc11p, a10=>pc10p, a9=>pc9p, a8=>pc8p, a7=>pc7p, a6=>pc6p);

  iwr_1f12 : ic_74s374 port map(oenb_n => gnd, o0 => iwr47, i0 => aa15, i1 => aa14, o1 => iwr46, o2 => iwr45, i2 => aa13, i3 => aa12, o3 => iwr44, clk => clk2c, o4 => iwr43, i4 => aa11, i5 => aa10, o5 => iwr42, o6 => iwr41, i6 => aa9, i7 => aa8, o7 => iwr40);
  iwr_1f14 : ic_74s374 port map(oenb_n => gnd, o0 => iwr39, i0 => aa7, i1 => aa6, o1 => iwr38, o2 => iwr37, i2 => aa5, i3 => aa4, o3 => iwr36, clk => clk2c, o4 => iwr35, i4 => aa3, i5 => aa2, o5 => iwr34, o6 => iwr33, i6 => aa1, i7 => aa0, o7 => iwr32);
  iwr_4b01 : ic_74s374 port map(oenb_n => gnd, o0 => iwr15, i0 => m15, i1 => m14, o1 => iwr14, o2 => iwr13, i2 => m13, i3 => m12, o3 => iwr12, clk => clk4c, o4 => iwr11, i4 => m11, i5 => m10, o5 => iwr10, o6 => iwr9, i6 => m9, i7 => m8, o7 => iwr8);
  iwr_4b06 : ic_74s374 port map(oenb_n => gnd, o0 => iwr7, i0 => m7, i1 => m6, o1 => iwr6, o2 => iwr5, i2 => m5, i3 => m4, o3 => iwr4, clk => clk4c, o4 => iwr3, i4 => m3, i5 => m2, o5 => iwr2, o6 => iwr1, i6 => m1, i7 => m0, o7 => iwr0);
  iwr_4c04 : ic_74s374 port map(oenb_n => gnd, o0 => iwr31, i0 => m31, i1 => m30, o1 => iwr30, o2 => iwr29, i2 => m29, i3 => m28, o3 => iwr28, clk => clk4c, o4 => iwr27, i4 => m27, i5 => m26, o5 => iwr26, o6 => iwr25, i6 => m25, i7 => m24, o7 => iwr24);
  iwr_4c05 : ic_74s374 port map(oenb_n => gnd, o0 => iwr23, i0 => m23, i1 => m22, o1 => iwr22, o2 => iwr21, i2 => m21, i3 => m20, o3 => iwr20, clk => clk4c, o4 => iwr19, i4 => m19, i5 => m18, o5 => iwr18, o6 => iwr17, i6 => m17, i7 => m16, o7 => iwr16);

  pctl_1a16 : ic_74ls244 port map(aenb_n => \-promenable\, ain0 => gnd, bout3 => nc29, ain1 => nc30, bout2 => nc31, ain2 => nc32, bout1 => nc33, ain3 => nc34, bout0 => nc35, bin0 => nc36, aout3 => nc37, bin1 => nc38, aout2 => nc39, bin2 => nc40, aout1 => nc41, bin3 => nc42, aout0 => i46, benb_n => hi2);
  pctl_1c17 : ic_74s04 port map(g1a      => pc0, g1q_n => \-prompc0\, g2a => pc1, g2q_n => \-prompc1\, g3a=>pc2, g3q_n=>\-prompc2\, g4q=>\-prompc3\, g4a=>pc3, g5q_n=>\-prompc4\, g5a=>pc4, g6q_n=>nc45, g6a=>nc46);
  pctl_1c18 : ic_74s32 port map(g1a      => \-promenable\, g1b => pc9, g1y => \-promce0\, g2a=>\-prompc9\, g2b=>\-promenable\, g2y=>\-promce1\, g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  pctl_1c19 : ic_74s20 port map(g1a      => \bottom.1k\, g1b => \-idebug\, g1c=>\-promdisabled\, g1d=>\-iwriteda\, g1y_n=>\-promenable\, g2a=>'0', g2b=>'0', g2c=>'0', g2d=>'0');
  pctl_1d18 : ic_74s260 port map(i1      => gnd, i2 => pc13, i3 => pc12, o1 => \bottom.1k\, i4 => pc11, i5 => pc10);
  pctl_1d19 : ic_74s04 port map(g1a      => pc5, g1q_n => \-prompc5\, g2a => pc6, g2q_n => \-prompc6\, g3a=>pc7, g3q_n=>\-prompc7\, g4q=>\-prompc8\, g4a=>pc8, g5q_n=>\-prompc9\, g5a=>pc9, g6q_n=>nc43, g6a=>nc44);
  pctl_1e16 : ic_74s20 port map(g1a      => \-ape\, g1b => \-pdlpe\, g1c=>\-spe\, g1d=>\-mpe\, g1y_n=>tilt1, g2y_n=>tilt0, g2a=>hi2, g2b=>\-mempe\, g2c=>\-v1pe\, g2d=>\-v0pe\);
  pctl_1f10 : ic_74s04 port map(g3a      => \-promenable\, g3q_n => promenable, g5q_n => dpe, g5a => \-dpe\, g6q_n=>ipe, g6a=>\-ipe\, g1a=>'0', g2a=>'0', g4a=>'0');
  pctl_1f16 : ic_til309 port map(l2      => nc4, l4 => nc5, l8 => nc6, l1 => nc7, latch => gnd, i4 => pc2, i8 => gnd, i2 => pc1, blank_n => hi2, dp => tilt1, test_n => hi2, ldp => nc8, i1 => pc0);
  pctl_1f17 : ic_til309 port map(l2      => nc9, l4 => nc10, l8 => nc11, l1 => nc12, latch => gnd, i4 => pc5, i8 => gnd, i2 => pc4, blank_n => hi2, dp => tilt0, test_n => hi2, ldp => nc13, i1 => pc3);
  pctl_1f18 : ic_til309 port map(l2      => nc14, l4 => nc15, l8 => nc16, l1 => nc17, latch => gnd, i4 => pc8, i8 => gnd, i2 => pc7, blank_n => hi2, dp => dpe, test_n => hi2, ldp => nc18, i1 => pc6);
  pctl_1f19 : ic_til309 port map(l2      => nc19, l4 => nc20, l8 => nc21, l1 => nc22, latch => gnd, i4 => pc11, i8 => gnd, i2 => pc10, blank_n => hi2, dp => ipe, test_n => hi2, ldp => nc23, i1 => pc9);
  pctl_1f20 : ic_til309 port map(l2      => nc24, l4 => nc25, l8 => nc26, l1 => nc27, latch => gnd, i4 => gnd, i8 => gnd, i2 => pc13, blank_n => hi2, dp => promenable, test_n => hi2, ldp => nc28, i1 => pc12);

  prom0_1b17 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i32, d1=>i33, d2=>i34, d3=>i35, d4=>i36, d5=>i37, d6=>i38, d7=>i39, ce_n=>\-promce0\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom0_1b19 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i40, d1=>i41, d2=>i42, d3=>i43, d4=>i44, d5=>i45, d6=>i47, d7=>i48, ce_n=>\-promce0\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom0_1c20 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i24, d1=>i25, d2=>i26, d3=>i27, d4=>i28, d5=>i29, d6=>i30, d7=>i31, ce_n=>\-promce0\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom0_1d16 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i16, d1=>i17, d2=>i18, d3=>i19, d4=>i20, d5=>i21, d6=>i22, d7=>i23, ce_n=>\-promce0\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom0_1e17 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i0, d1=>i1, d2=>i2, d3=>i3, d4=>i4, d5=>i5, d6=>i6, d7=>i7, ce_n=>\-promce0\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom0_1e19 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i8, d1=>i9, d2=>i10, d3=>i11, d4=>i12, d5=>i13, d6=>i14, d7=>i15, ce_n=>\-promce0\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);

  prom1_1b16 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i24, d1=>i25, d2=>i26, d3=>i27, d4=>i28, d5=>i29, d6=>i30, d7=>i31, ce_n=>\-promce1\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom1_1b18 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i32, d1=>i33, d2=>i34, d3=>i35, d4=>i36, d5=>i37, d6=>i38, d7=>i39, ce_n=>\-promce1\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom1_1b20 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i40, d1=>i41, d2=>i42, d3=>i43, d4=>i44, d5=>i45, d6=>i47, d7=>i48, ce_n=>\-promce1\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom1_1d17 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i16, d1=>i17, d2=>i18, d3=>i19, d4=>i20, d5=>i21, d6=>i22, d7=>i23, ce_n=>\-promce1\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom1_1e18 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i0, d1=>i1, d2=>i2, d3=>i3, d4=>i4, d5=>i5, d6=>i6, d7=>i7, ce_n=>\-promce1\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);
  prom1_1e20 : ic_74s472 port map(a0 => \-prompc0\, a1 => \-prompc1\, a2=>\-prompc2\, a3=>\-prompc3\, a4=>\-prompc4\, d0=>i8, d1=>i9, d2=>i10, d3=>i11, d4=>i12, d5=>i13, d6=>i14, d7=>i15, ce_n=>\-promce1\, a5=>\-prompc5\, a6=>\-prompc6\, a7=>\-prompc7\, a8=>\-prompc8\);

  debug_1e11 : ic_74s374 port map(oenb_n => \-idebug\, o0 => i39, i0 => spy7, i1 => spy6, o1 => i38, o2 => i37, i2 => spy5, i3 => spy4, o3 => i36, clk => \-lddbirh\, o4=>i35, i4=>spy3, i5=>spy2, o5=>i34, o6=>i33, i6=>spy1, i7=>spy0, o7=>i32);
  debug_1e12 : ic_74s374 port map(oenb_n => \-idebug\, o0 => i31, i0 => spy15, i1 => spy14, o1 => i30, o2 => i29, i2 => spy13, i3 => spy12, o3 => i28, clk => \-lddbirm\, o4=>i27, i4=>spy11, i5=>spy10, o5=>i26, o6=>i25, i6=>spy9, i7=>spy8, o7=>i24);
  debug_1e13 : ic_74s374 port map(oenb_n => \-idebug\, o0 => i23, i0 => spy7, i1 => spy6, o1 => i22, o2 => i21, i2 => spy5, i3 => spy4, o3 => i20, clk => \-lddbirm\, o4=>i19, i4=>spy3, i5=>spy2, o5=>i18, o6=>i17, i6=>spy1, i7=>spy0, o7=>i16);
  debug_1e14 : ic_74s374 port map(oenb_n => \-idebug\, o0 => i15, i0 => spy15, i1 => spy14, o1 => i14, o2 => i13, i2 => spy13, i3 => spy12, o3 => i12, clk => \-lddbirl\, o4=>i11, i4=>spy11, i5=>spy10, o5=>i10, o6=>i9, i6=>spy9, i7=>spy8, o7=>i8);
  debug_1e15 : ic_74s374 port map(oenb_n => \-idebug\, o0 => i7, i0 => spy7, i1 => spy6, o1 => i6, o2 => i5, i2 => spy5, i3 => spy4, o3 => i4, clk => \-lddbirl\, o4=>i3, i4=>spy3, i5=>spy2, o5=>i2, o6=>i1, i6=>spy1, i7=>spy0, o7=>i0);
  debug_1f15 : ic_74s374 port map(oenb_n => \-idebug\, o0 => i47, i0 => spy15, i1 => spy14, o1 => i46, o2 => i45, i2 => spy13, i3 => spy12, o3 => i44, clk => \-lddbirh\, o4=>i43, i4=>spy11, i5=>spy10, o5=>i42, o6=>i41, i6=>spy9, i7=>spy8, o7=>i40);

  --- Microinstrction Modification and Main Instruction Register

  ior_3c06 : ic_74s32 port map(g1a => i12, g1b => ob12, g1y => iob12, g2a => i13, g2b => ob13, g2y => iob13, g3y => iob14, g3a => i14, g3b => ob14, g4y => iob15, g4a => i15, g4b => ob15);
  ior_3c07 : ic_74s32 port map(g1a => i8, g1b => ob8, g1y => iob8, g2a => i9, g2b => ob9, g2y => iob9, g3y => iob10, g3a => i10, g3b => ob10, g4y => iob11, g4a => i11, g4b => ob11);
  ior_3c08 : ic_74s32 port map(g1a => i4, g1b => ob4, g1y => iob4, g2a => i5, g2b => ob5, g2y => iob5, g3y => iob6, g3a => i6, g3b => ob6, g4y => iob7, g4a => i7, g4b => ob7);
  ior_3c09 : ic_74s32 port map(g1a => i0, g1b => ob0, g1y => iob0, g2a => i1, g2b => ob1, g2y => iob1, g3y => iob2, g3a => i2, g3b => ob2, g4y => iob3, g4a => i3, g4b => ob3);
  ior_3c16 : ic_74s32 port map(g1a => i20, g1b => ob20, g1y => iob20, g2a => i21, g2b => ob21, g2y => iob21, g3y => iob22, g3a => i22, g3b => ob22, g4y => iob23, g4a => i23, g4b => ob23);
  ior_3c18 : ic_74s32 port map(g1a => i16, g1b => ob16, g1y => iob16, g2a => i17, g2b => ob17, g2y => iob17, g3y => iob18, g3a => i18, g3b => ob18, g4y => iob19, g4a => i19, g4b => ob19);
  ior_3d08 : ic_74s32 port map(g1a => i44, g1b => ob18, g1y => iob44, g2a => i45, g2b => ob19, g2y => iob45, g3y => iob46, g3a => i46, g3b => ob20, g4y => iob47, g4a => i47, g4b => ob21);
  ior_3d09 : ic_74s32 port map(g1a => i40, g1b => ob14, g1y => iob40, g2a => i41, g2b => ob15, g2y => iob41, g3y => iob42, g3a => i42, g3b => ob16, g4y => iob43, g4a => i43, g4b => ob17);
  ior_3d10 : ic_74s32 port map(g1a => i36, g1b => ob10, g1y => iob36, g2a => i37, g2b => ob11, g2y => iob37, g3y => iob38, g3a => i38, g3b => ob12, g4y => iob39, g4a => i39, g4b => ob13);
  ior_3d13 : ic_74s32 port map(g1a => i32, g1b => ob6, g1y => iob32, g2a => i33, g2b => ob7, g2y => iob33, g3y => iob34, g3a => i34, g3b => ob8, g4y => iob35, g4a => i35, g4b => ob9);
  ior_3d14 : ic_74s32 port map(g1a => i28, g1b => ob2, g1y => iob28, g2a => i29, g2b => ob3, g2y => iob29, g3y => iob30, g3a => i30, g3b => ob4, g4y => iob31, g4a => i31, g4b => ob5);
  ior_3d15 : ic_74s32 port map(g1a => i24, g1b => ob24, g1y => iob24, g2a => i25, g2b => ob25, g2y => iob25, g3y => iob26, g3a => i26, g3b => ob0, g4y => iob27, g4a => i27, g4b => ob1);

  ireg_3c01 : ic_25s09 port map(sel => \-destimod0\, aq => ir15, a0 => iob15, a1 => i15, b1 => i14, b0 => iob14, bq => ir14, clk => clk3a, cq => ir13, c0 => iob13, c1 => i13, d1 => i12, d0 => iob12, dq => ir12);
  ireg_3c02 : ic_25s09 port map(sel => \-destimod0\, aq => ir11, a0 => iob11, a1 => i11, b1 => i10, b0 => iob10, bq => ir10, clk => clk3a, cq => ir9, c0 => iob9, c1 => i9, d1 => i8, d0 => iob8, dq => ir8);
  ireg_3c03 : ic_25s09 port map(sel => \-destimod0\, aq => ir7, a0 => iob7, a1 => i7, b1 => i6, b0 => iob6, bq => ir6, clk => clk3a, cq => ir5, c0 => iob5, c1 => i5, d1 => i4, d0 => iob4, dq => ir4);
  ireg_3c04 : ic_25s09 port map(sel => \-destimod0\, aq => ir3, a0 => iob3, a1 => i3, b1 => i2, b0 => iob2, bq => ir2, clk => clk3a, cq => ir1, c0 => iob1, c1 => i1, d1 => i0, d0 => iob0, dq => ir0);
  ireg_3c17 : ic_25s09 port map(sel => \-destimod0\, aq => ir23, a0 => iob23, a1 => i23, b1 => i22, b0 => iob22, bq => ir22, clk => clk3b, cq => ir21, c0 => iob21, c1 => i21, d1 => i20, d0 => iob20, dq => ir20);
  ireg_3c19 : ic_25s09 port map(sel => \-destimod0\, aq => ir19, a0 => iob19, a1 => i19, b1 => i18, b0 => iob18, bq => ir18, clk => clk3b, cq => ir17, c0 => iob17, c1 => i17, d1 => i16, d0 => iob16, dq => ir16);
  ireg_3d06 : ic_25s09 port map(sel => \-destimod1\, aq => nc371, a0 => nc372, a1 => nc373, b1 => i48, b0 => gnd, bq => ir48, clk => clk3a, cq => ir47, c0 => iob47, c1 => i47, d1 => i46, d0 => iob46, dq => ir46);
  ireg_3d07 : ic_25s09 port map(sel => \-destimod1\, aq => ir45, a0 => iob45, a1 => i45, b1 => i44, b0 => iob44, bq => ir44, clk => clk3a, cq => ir43, c0 => iob43, c1 => i43, d1 => i42, d0 => iob42, dq => ir42);
  ireg_3d16 : ic_25s09 port map(sel => \-destimod1\, aq => ir41, a0 => iob41, a1 => i41, b1 => i40, b0 => iob40, bq => ir40, clk => clk3b, cq => ir39, c0 => iob39, c1 => i39, d1 => i38, d0 => iob38, dq => ir38);
  ireg_3d17 : ic_25s09 port map(sel => \-destimod1\, aq => ir37, a0 => iob37, a1 => i37, b1 => i36, b0 => iob36, bq => ir36, clk => clk3b, cq => ir35, c0 => iob35, c1 => i35, d1 => i34, d0 => iob34, dq => ir34);
  ireg_3d18 : ic_25s09 port map(sel => \-destimod1\, aq => ir33, a0 => iob33, a1 => i33, b1 => i32, b0 => iob32, bq => ir32, clk => clk3b, cq => ir31, c0 => iob31, c1 => i31, d1 => i30, d0 => iob30, dq => ir30);
  ireg_3d19 : ic_25s09 port map(sel => \-destimod1\, aq => ir29, a0 => iob29, a1 => i29, b1 => i28, b0 => iob28, bq => ir28, clk => clk3b, cq => ir27, c0 => iob27, c1 => i27, d1 => i26, d0 => iob26, dq => ir26);
  ireg_3d20 : ic_25s09 port map(sel => \-destimod0\, aq => nc374, a0 => nc375, a1 => nc376, b1 => nc377, b0 => nc378, bq => nc379, clk => clk3b, cq => ir25, c0 => iob25, c1 => i25, d1 => i24, d0 => iob24, dq => ir24);

  --- IR Decoding

  source_3d02 : ic_74s00 port map(g2b => \-iralu\, g2a => \-irbyte\, g2q_n=>dest, g3q_n=>\-destmem\, g3b=>ir23, g3a=>destm, g4q_n=>\-specalu\, g4a=>ir8, g4b=>iralu, g1b=>'0', g1a=>'0');
  source_3d03 : ic_74s04 port map(g1a => ir22, g1q_n => \-ir22\, g2a => ir25, g2q_n => \-ir25\, g3a=>nc198, g3q_n=>nc199, g4q=>irdisp, g4a=>\-irdisp\, g5q_n=>irjump, g5a=>\-irjump\, g6q_n=>iralu, g6a=>\-iralu\);
  source_3d04 : ic_74s139 port map(g1 => \-specalu\, a1 => ir3, b1 => ir4, g1y0 => \-mul\, g1y1=>\-div\, g1y2=>nc196, g1y3=>nc197, b2=>'0', a2=>'0', g2=>'0');
  source_3d05 : ic_74s139 port map(g1 => nop, a1 => ir43, b1 => ir44, g1y0 => \-iralu\, g1y1 => \-irjump\, g1y2=>\-irdisp\, g1y3=>\-irbyte\, g2y3=>\-funct3\, g2y2=>\-funct2\, g2y1=>\-funct1\, g2y0=>\-funct0\, b2=>ir11, a2=>ir10, g2=>nop);
  source_3d11 : ic_74s138 port map(a  => ir19, b => ir20, c => ir21, g2a => ir22, g2b => ir23, g1 => destm, y7 => nc200, y6 => nc201, y5 => nc202, y4 => nc203, y3 => nc204, y2 => \-destintctl\, y1 => \-destlc\, y0=>nc205);
  source_3d12 : ic_74s138 port map(a  => ir19, b => ir20, c => ir21, g2a => \-ir22\, g2b => ir23, g1 => destm, y7 => \-destimod1\, y6=>\-destimod0\, y5=>\-destspc\, y4=>\-destpdlp\, y3=>\-destpdlx\, y2=>\-destpdl(x)\, y1=>\-destpdl(p)\, y0=>\-destpdltop\);
  source_3d21 : ic_74s08 port map(g4q => destm, g4a => \-ir25\, g4b => dest, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3a => '0', g3b => '0');
  source_3d22 : ic_74s138 port map(a  => ir26, b => ir27, c => ir28, g2a => \-ir31\, g2b => ir29, g1 => hi5, y7 => \-srcq\, y6=>\-srcopc\, y5=>\-srcpdltop\, y4=>\-srcpdlpop\, y3=>\-srcpdlidx\, y2=>\-srcpdlptr\, y1=>\-srcspc\, y0=>\-srcdc\);
  source_3d23 : ic_74s138 port map(a  => ir26, b => ir27, c => ir28, g2a => \-ir31\, g2b => gnd, g1 => ir29, y7 => nc206, y6 => nc207, y5 => nc208, y4 => \-srcspcpop\, y3=>\-srclc\, y2=>\-srcmd\, y1=>\-srcmap\, y0=>\-srcvma\);
  source_3e05 : ic_74s08 port map(g2b => \destimod0_l\, g2a => \iwrited_l\, g2q=>internal18, g1b=>'0', g1a=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  source_3e09 : ic_74s32 port map(g2a => \-destmem\, g2b => \-ir22\, g2y=>\-destmdr\, g3y=>\-destvma\, g3a=>ir22, g3b=>\-destmem\, g1a=>'0', g1b=>'0', g4a=>'0', g4b=>'0');
  source_4d10 : ic_74s10 port map(g2a => internal18, g2b => \-destimod1\, g2c => \-idebug\, g2y_n=>imod, g1a=>'0', g1b=>'0', g3a=>'0', g3b=>'0', g3c=>'0', g1c=>'0');

  --- A Memory

  actl_3a06 : ic_74s258 port map(sel   => clk3e, d0 => wadr0, d1 => ir32, dy => \-aadr0b\, c0 => wadr1, c1 => ir33, cy => \-aadr1b\, by=>\-aadr2b\, b1=>ir34, b0=>wadr2, ay=>\-aadr3b\, a1=>ir35, a0=>wadr3, enb_n=>gnd);
  actl_3a12 : ic_74s258 port map(sel   => clk3d, d0 => wadr4, d1 => ir36, dy => \-aadr4b\, c0 => wadr5, c1 => ir37, cy => \-aadr5b\, by=>\-aadr6b\, b1=>ir38, b0=>wadr6, ay=>\-aadr7b\, a1=>ir39, a0=>wadr7, enb_n=>gnd);
  actl_3a16 : ic_74s258 port map(sel   => clk3d, d0 => wadr0, d1 => ir32, dy => \-aadr0a\, c0 => wadr1, c1 => ir33, cy => \-aadr1a\, by=>\-aadr2a\, b1=>ir34, b0=>wadr2, ay=>\-aadr3a\, a1=>ir35, a0=>wadr3, enb_n=>gnd);
  actl_3a21 : ic_74s258 port map(sel   => clk3d, d0 => wadr4, d1 => ir36, dy => \-aadr4a\, c0 => wadr5, c1 => ir37, cy => \-aadr5a\, by=>\-aadr6a\, b1=>ir38, b0=>wadr6, ay=>\-aadr7a\, a1=>ir39, a0=>wadr7, enb_n=>gnd);
  actl_3b15 : ic_74s258 port map(sel   => clk3d, d0 => wadr8, d1 => ir40, dy => \-aadr8a\, c0 => wadr9, c1 => ir41, cy => \-aadr9a\, by=>\-aadr8b\, b1=>ir40, b0=>wadr8, ay=>\-aadr9b\, a1=>ir41, a0=>wadr9, enb_n=>gnd);
  actl_3b16 : ic_74s00 port map(g1b    => apass1, g1a => apass2, g1q_n => \-apass\, g2b => \-apass\, g2a=>tse3a, g2q_n=>\-amemenb\, g3b=>'0', g3a=>'0', g4a=>'0', g4b=>'0');
  actl_3b21 : ic_93s46 port map(a0     => ir32, b0 => wadr0, a1 => ir33, b1 => wadr1, a2 => ir34, b2 => wadr2, enb => hi3, eq => apass1, a3 => ir35, b3 => wadr3, a4 => ir36, b4 => wadr4, a5 => ir37, b5 => wadr5);
  actl_3b26 : ic_74s174 port map(clr_n => \-reset\, q1 => wadr0, d1 => ir14, d2 => ir15, q2 => wadr1, d3 => ir16, q3 => wadr2, clk => clk3d, q4 => wadr3, d4 => ir17, q5 => destmd, d5 => destm, d6 => dest, q6 => destd);
  actl_3b27 : ic_93s46 port map(a0     => ir38, b0 => wadr6, a1 => ir39, b1 => wadr7, a2 => ir40, b2 => wadr8, enb => hi3, eq => apass2, a3 => ir41, b3 => wadr9, a4 => hi3, b4 => destd, a5 => gnd, b5 => gnd);
  actl_3b28 : ic_25s09 port map(sel    => destm, aq => wadr7, a0 => ir21, a1 => gnd, b1 => gnd, b0 => ir20, bq => wadr6, clk => clk3d, cq => wadr5, c0 => ir19, c1 => gnd, d1 => ir18, d0 => ir18, dq => wadr4);
  actl_3b29 : ic_25s09 port map(sel    => destm, aq => nc489, a0 => nc490, a1 => nc491, b1 => nc492, b0 => nc493, bq => nc494, clk => clk3d, cq => wadr9, c0 => ir23, c1 => gnd, d1 => gnd, d0 => ir22, dq => wadr8);
  actl_3b30 : ic_74s37 port map(g1a    => wp3a, g1b => destd, g1y => \-awpa\, g2a => wp3a, g2b => destd, g2y => \-awpb\, g3y=>\-awpc\, g3a=>destd, g3b=>wp3a, g4a=>'0', g4b=>'0');
  actl_4b11 : ic_74s11 port map(g2a    => apass1, g2b => apass2, g2c => tse4a, g2y_n => apassenb, g1a => '0', g1b => '0', g3a => '0', g3b => '0', g3c => '0', g1c => '0');
  actl_4b14 : ic_74s10 port map(g3y_n  => \-apassenb\, g3a => tse4a, g3b => apass2, g3c => apass1, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g2c => '0', g1c => '0');

  amem0_3a07 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem22, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l22);
  amem0_3a08 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem20, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l20);
  amem0_3a09 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem18, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l18);
  amem0_3a10 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem16, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l16);
  amem0_3a11 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem23, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l23);
  amem0_3a13 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem21, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l21);
  amem0_3a14 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem19, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l19);
  amem0_3a15 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem17, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l17);
  amem0_3b06 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amemparity, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>lparity);
  amem0_3b07 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem30, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l30);
  amem0_3b08 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem28, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l28);
  amem0_3b09 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem26, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l26);
  amem0_3b10 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem24, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l24);
  amem0_3b11 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem31, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l31);
  amem0_3b12 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem29, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l29);
  amem0_3b13 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem27, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l27);
  amem0_3b14 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0b\, a1 => \-aadr1b\, a2=>\-aadr2b\, a3=>\-aadr3b\, a4=>\-aadr4b\, do=>amem25, a5=>\-aadr5b\, a6=>\-aadr6b\, a7=>\-aadr7b\, a8=>\-aadr8b\, a9=>\-aadr9b\, we_n=>\-awpa\, di=>l25);

  amem1_3a17 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem6, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l6);
  amem1_3a18 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem4, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l4);
  amem1_3a19 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem2, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l2);
  amem1_3a20 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem0, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l0);
  amem1_3a22 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem7, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l7);
  amem1_3a23 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem5, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l5);
  amem1_3a24 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem3, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l3);
  amem1_3a25 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem1, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l1);
  amem1_3b17 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem14, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpb\, di=>l14);
  amem1_3b18 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem12, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpb\, di=>l12);
  amem1_3b19 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem10, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l10);
  amem1_3b20 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem8, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l8);
  amem1_3b22 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem15, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpb\, di=>l15);
  amem1_3b23 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem13, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpb\, di=>l13);
  amem1_3b24 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem11, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpb\, di=>l11);
  amem1_3b25 : ic_93425a port map(ce_n => gnd, a0 => \-aadr0a\, a1 => \-aadr1a\, a2=>\-aadr2a\, a3=>\-aadr3a\, a4=>\-aadr4a\, do=>amem9, a5=>\-aadr5a\, a6=>\-aadr6a\, a7=>\-aadr7a\, a8=>\-aadr8a\, a9=>\-aadr9a\, we_n=>\-awpc\, di=>l9);

  alatch_3a01 : ic_74s373 port map(oenb_n => \-amemenb\, o0 => a23, i0 => amem23, i1 => amem22, o1 => a22, o2 => a21, i2 => amem21, i3 => amem20, o3 => a20, hold_n => clk3e, o4 => a19, i4 => amem19, i5 => amem18, o5 => a18, o6 => a17, i6 => amem17, i7 => amem16, o7 => a16);
  alatch_3a02 : ic_74s241 port map(aenb_n => \-apassenb\, ain0 => l15, bout3 => a8, ain1 => l14, bout2 => a9, ain2 => l13, bout1 => a10, ain3 => l12, bout0 => a11, bin0 => l11, aout3 => a12, bin1 => l10, aout2 => a13, bin2 => l9, aout1 => a14, bin3 => l8, aout0 => a15, benb => apassenb);
  alatch_3a03 : ic_74s373 port map(oenb_n => \-amemenb\, o0 => a15, i0 => amem15, i1 => amem14, o1 => a14, o2 => a13, i2 => amem13, i3 => amem12, o3 => a12, hold_n => clk3e, o4 => a11, i4 => amem11, i5 => amem10, o5 => a10, o6 => a9, i6 => amem9, i7 => amem8, o7 => a8);
  alatch_3a04 : ic_74s241 port map(aenb_n => \-apassenb\, ain0 => l7, bout3 => a0, ain1 => l6, bout2 => a1, ain2 => l5, bout1 => a2, ain3 => l4, bout0 => a3, bin0 => l3, aout3 => a4, bin1 => l2, aout2 => a5, bin2 => l1, aout1 => a6, bin3 => l0, aout0 => a7, benb => apassenb);
  alatch_3a05 : ic_74s373 port map(oenb_n => \-amemenb\, o0 => a7, i0 => amem7, i1 => amem6, o1 => a6, o2 => a5, i2 => amem5, i3 => amem4, o3 => a4, hold_n => clk3e, o4 => a3, i4 => amem3, i5 => amem2, o5 => a2, o6 => a1, i6 => amem1, i7 => amem0, o7 => a0);
  alatch_3b01 : ic_74s241 port map(aenb_n => hi5, ain0 => nc465, bout3 => a31b, ain1 => nc466, bout2 => aparity, ain2 => nc467, bout1 => nc468, ain3 => nc469, bout0 => nc470, bin0 => nc471, aout3 => nc472, bin1 => nc473, aout2 => nc474, bin2 => lparity, aout1 => nc475, bin3 => l31, aout0 => nc476, benb => apassenb);
  alatch_3b02 : ic_74s373 port map(oenb_n => \-amemenb\, o0 => nc477, i0 => nc478, i1 => nc479, o1 => nc480, o2 => nc481, i2 => nc482, i3 => nc483, o3 => nc484, hold_n => clk3e, o4 => nc485, i4 => nc486, i5 => nc487, o5 => nc488, o6 => aparity, i6 => amemparity, i7 => amem31, o7 => a31b);
  alatch_3b03 : ic_74s241 port map(aenb_n => \-apassenb\, ain0 => l31, bout3 => a24, ain1 => l30, bout2 => a25, ain2 => l29, bout1 => a26, ain3 => l28, bout0 => a27, bin0 => l27, aout3 => a28, bin1 => l26, aout2 => a29, bin2 => l25, aout1 => a30, bin3 => l24, aout0 => a31a, benb => apassenb);
  alatch_3b04 : ic_74s373 port map(oenb_n => \-amemenb\, o0 => a31a, i0 => amem31, i1 => amem30, o1 => a30, o2 => a29, i2 => amem29, i3 => amem28, o3 => a28, hold_n => clk3e, o4 => a27, i4 => amem27, i5 => amem26, o5 => a26, o6 => a25, i6 => amem25, i7 => amem24, o7 => a24);
  alatch_3b05 : ic_74s241 port map(aenb_n => \-apassenb\, ain0 => l23, bout3 => a16, ain1 => l22, bout2 => a17, ain2 => l21, bout1 => a18, ain3 => l20, bout0 => a19, bin0 => l19, aout3 => a20, bin1 => l18, aout2 => a21, bin2 => l17, aout1 => a22, bin3 => l16, aout0 => a23, benb => apassenb);

  apar_3a28 : ic_93s48 port map(i6  => a26, i5 => a27, i4 => a28, i3 => a29, i2 => a30, i1 => a31b, i0 => aparity, po => aparok, pe => nc432, i11 => aparl, i10 => aparm, i9 => gnd, i8 => a24, i7 => a25);
  apar_3a29 : ic_93s48 port map(i6  => a17, i5 => a18, i4 => a19, i3 => a20, i2 => a21, i1 => a22, i0 => a23, po => aparm, pe => nc433, i11 => a12, i10 => a13, i9 => a14, i8 => a15, i7 => a16);
  apar_3a30 : ic_93s48 port map(i6  => a5, i5 => a6, i4 => a7, i3 => a8, i2 => a9, i1 => a10, i0 => a11, po => aparl, pe => nc434, i11 => a0, i10 => a1, i9 => a2, i8 => a3, i7 => a4);
  apar_4a12 : ic_93s48 port map(i6  => m17, i5 => m18, i4 => m19, i3 => m20, i2 => m21, i1 => m22, i0 => m23, po => mparm, pe => nc436, i11 => m12, i10 => m13, i9 => m14, i8 => m15, i7 => m16);
  apar_4a14 : ic_93s48 port map(i6  => m5, i5 => m6, i4 => m7, i3 => m8, i2 => m9, i1 => m10, i0 => m11, po => mparl, pe => nc435, i11 => m0, i10 => m1, i9 => m2, i8 => m3, i7 => m4);
  apar_4a17 : ic_74s00 port map(g1b => mpareven, g1a => srcm, g1q_n => mmemparok, g2b => mpareven, g2a => pdlenb, g2q_n => pdlparok, g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  apar_4b15 : ic_93s48 port map(i6  => m26, i5 => m27, i4 => m28, i3 => m29, i2 => m30, i1 => m31, i0 => mparity, po => mparodd, pe => mpareven, i11 => mparl, i10 => mparm, i9 => gnd, i8 => m24, i7 => m25);

  --- M Memory

  mctl_4a16 : ic_74s258 port map(sel => clk4e, d0 => wadr4, d1 => ir30, dy => \-madr4a\, c0 => nc335, c1 => nc336, cy => nc337, by => nc338, b1 => nc339, b0 => nc340, ay => \-madr4b\, a1=>ir30, a0=>wadr4, enb_n=>gnd);
  mctl_4a18 : ic_74s258 port map(sel => clk4e, d0 => wadr0, d1 => ir26, dy => \-madr0b\, c0 => wadr1, c1 => ir27, cy => \-madr1b\, by=>\-madr2b\, b1=>ir28, b0=>wadr2, ay=>\-madr3b\, a1=>ir29, a0=>wadr3, enb_n=>gnd);
  mctl_4a19 : ic_res20 port map(r2   => nc334, r3 => mmem15, r4 => mmem14, r5 => mmem13, r6 => mmem12, r7 => mmem11, r8 => mmem10, r9 => mmem9, r11 => mmem8, r12 => mmem7, r13 => mmem6, r14 => mmem5, r15 => mmem4, r16 => mmem3, r17 => mmem2, r18 => mmem1, r19 => mmem0, r10 => '0');
  mctl_4b11 : ic_74s11 port map(g1a  => mpass, g1b => tse4a, g3y_n => srcm, g3a => hi2, g3b => \-ir31\, g3c => \-mpass\, g1y_n=>mpassl, g1c=>\-ir31\, g2a=>'0', g2b=>'0', g2c=>'0');
  mctl_4b12 : ic_74s04 port map(g1a  => mpass, g1q_n => \-mpass\, g2a => '0', g3a => '0', g4a => '0', g5a => '0', g6a => '0');
  mctl_4b14 : ic_74s10 port map(g1a  => mpass, g1b => tse4a, g2a => tse4a, g2b => \-ir31\, g2c => \-mpass\, g2y_n=>\-mpassm\, g1y_n=>\-mpassl\, g1c=>\-ir31\, g3a=>'0', g3b=>'0', g3c=>'0');
  mctl_4b18 : ic_93s46 port map(a0   => ir26, b0 => wadr0, a1 => ir27, b1 => wadr1, a2 => ir28, b2 => wadr2, enb => hi2, eq => mpass, a3 => ir29, b3 => wadr3, a4 => ir30, b4 => wadr4, a5 => hi2, b5 => destmd);
  mctl_4b19 : ic_74s258 port map(sel => clk4e, d0 => wadr0, d1 => ir26, dy => \-madr0a\, c0 => wadr1, c1 => ir27, cy => \-madr1a\, by=>\-madr2a\, b1=>ir28, b0=>wadr2, ay=>\-madr3a\, a1=>ir29, a0=>wadr3, enb_n=>gnd);
  mctl_4b20 : ic_res20 port map(r2   => mmemparity, r3 => mmem31, r4 => mmem30, r5 => mmem29, r6 => mmem28, r7 => mmem27, r8 => mmem26, r9 => mmem25, r11 => mmem24, r12 => mmem23, r13 => mmem22, r14 => mmem21, r15 => mmem20, r16 => mmem19, r17 => mmem18, r18 => mmem17, r19 => mmem16, r10 => '0');
  mctl_4b22 : ic_74s37 port map(g1a  => destmd, g1b => wp4b, g1y => \-mwpa\, g2a => destmd, g2b => wp4b, g2y => \-mwpb\, g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');

  mmem_4a21 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l16, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem16, d1=>mmem17, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l17, we1_n=>gnd);
  mmem_4a22 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l12, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem12, d1=>mmem13, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l13, we1_n=>gnd);
  mmem_4a23 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l8, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem8, d1=>mmem9, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l9, we1_n=>gnd);
  mmem_4a24 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l4, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem4, d1=>mmem5, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l5, we1_n=>gnd);
  mmem_4a25 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l0, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem0, d1=>mmem1, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l1, we1_n=>gnd);
  mmem_4a26 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l18, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem18, d1=>mmem19, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l19, we1_n=>gnd);
  mmem_4a27 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l14, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem14, d1=>mmem15, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l15, we1_n=>gnd);
  mmem_4a28 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l10, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem10, d1=>mmem11, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l11, we1_n=>gnd);
  mmem_4a29 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l6, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem6, d1=>mmem7, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l7, we1_n=>gnd);
  mmem_4a30 : ic_82s21 port map(wclk_n => \-mwpb\, we0_n => gnd, i0 => l2, a4 => \-madr4b\, ce=>hi2, strobe=>hi2, d0=>mmem2, d1=>mmem3, a3=>\-madr3b\, a2=>\-madr2b\, a1=>\-madr1b\, a0=>\-madr0b\, i1=>l3, we1_n=>gnd);
  mmem_4b23 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l28, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem28, d1=>mmem29, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l29, we1_n=>gnd);
  mmem_4b24 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l24, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem24, d1=>mmem25, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l25, we1_n=>gnd);
  mmem_4b25 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l20, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem20, d1=>mmem21, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l21, we1_n=>gnd);
  mmem_4b27 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => lparity, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmemparity, d1=>nc291, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>nc292, we1_n=>nc293);
  mmem_4b28 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l30, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem30, d1=>mmem31, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l31, we1_n=>gnd);
  mmem_4b29 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l26, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem26, d1=>mmem27, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l27, we1_n=>gnd);
  mmem_4b30 : ic_82s21 port map(wclk_n => \-mwpa\, we0_n => gnd, i0 => l22, a4 => \-madr4a\, ce=>hi3, strobe=>hi3, d0=>mmem22, d1=>mmem23, a3=>\-madr3a\, a2=>\-madr2a\, a1=>\-madr1a\, a0=>\-madr0a\, i1=>l23, we1_n=>gnd);

  mlatch_4a01 : ic_74s373 port map(oenb_n => \-mpassm\, o0 => m23, i0 => mmem23, i1 => mmem22, o1 => m22, o2 => m21, i2 => mmem21, i3 => mmem20, o3 => m20, hold_n => clk4a, o4 => m19, i4 => mmem19, i5 => mmem18, o5 => m18, o6 => m17, i6 => mmem17, i7 => mmem16, o7 => m16);
  mlatch_4a03 : ic_74s373 port map(oenb_n => \-mpassm\, o0 => m15, i0 => mmem15, i1 => mmem14, o1 => m14, o2 => m13, i2 => mmem13, i3 => mmem12, o3 => m12, hold_n => clk4a, o4 => m11, i4 => mmem11, i5 => mmem10, o5 => m10, o6 => m9, i6 => mmem9, i7 => mmem8, o7 => m8);
  mlatch_4a05 : ic_74s373 port map(oenb_n => \-mpassm\, o0 => m7, i0 => mmem7, i1 => mmem6, o1 => m6, o2 => m5, i2 => mmem5, i3 => mmem4, o3 => m4, hold_n => clk4a, o4 => m3, i4 => mmem3, i5 => mmem2, o5 => m2, o6 => m1, i6 => mmem1, i7 => mmem0, o7 => m0);
  mlatch_4a06 : ic_74s241 port map(aenb_n => \-mpassl\, ain0 => l15, bout3 => mf8, ain1 => l14, bout2 => mf9, ain2 => l13, bout1 => mf10, ain3 => l12, bout0 => mf11, bin0 => l11, aout3 => mf12, bin1 => l10, aout2 => mf13, bin2 => l9, aout1 => mf14, bin3 => l8, aout0 => mf15, benb => mpassl);
  mlatch_4a08 : ic_74s241 port map(aenb_n => \-mpassl\, ain0 => l7, bout3 => mf0, ain1 => l6, bout2 => mf1, ain2 => l5, bout1 => mf2, ain3 => l4, bout0 => mf3, bin0 => l3, aout3 => mf4, bin1 => l2, aout2 => mf5, bin2 => l1, aout1 => mf6, bin3 => l0, aout0 => mf7, benb => mpassl);
  mlatch_4b02 : ic_74s373 port map(oenb_n => \-mpassm\, o0 => nc294, i0 => nc295, i1 => nc296, o1 => nc297, o2 => nc298, i2 => nc299, i3 => nc300, o3 => nc301, hold_n => clk4a, o4 => nc302, i4 => nc303, i5 => nc304, o5 => nc305, o6 => nc306, i6 => nc307, i7 => mmemparity, o7 => mparity);
  mlatch_4b04 : ic_74s373 port map(oenb_n => \-mpassm\, o0 => m31, i0 => mmem31, i1 => mmem30, o1 => m30, o2 => m29, i2 => mmem29, i3 => mmem28, o3 => m28, hold_n => clk4a, o4 => m27, i4 => mmem27, i5 => mmem26, o5 => m26, o6 => m25, i6 => mmem25, i7 => mmem24, o7 => m24);
  mlatch_4b07 : ic_74s241 port map(aenb_n => \-mpassl\, ain0 => l31, bout3 => mf24, ain1 => l30, bout2 => mf25, ain2 => l29, bout1 => mf26, ain3 => l28, bout0 => mf27, bin0 => l27, aout3 => mf28, bin1 => l26, aout2 => mf29, bin2 => l25, aout1 => mf30, bin3 => l24, aout0 => mf31, benb => mpassl);
  mlatch_4b09 : ic_74s241 port map(aenb_n => \-mpassl\, ain0 => l23, bout3 => mf16, ain1 => l22, bout2 => mf17, ain2 => l21, bout1 => mf18, ain3 => l20, bout0 => mf19, bin0 => l19, aout3 => mf20, bin1 => l18, aout2 => mf21, bin2 => l17, aout1 => mf22, bin3 => l16, aout0 => mf23, benb => mpassl);

  mf_1a18 : ic_74s00 port map(g1b     => tse1a, g1a => mfenb, g1q_n => \-mfdrive\, g2b => '0', g2a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  mf_1a21 : ic_74s241 port map(aenb_n => \-mfdrive\, ain0 => mf23, bout3 => m16, ain1 => mf22, bout2 => m17, ain2 => mf21, bout1 => m18, ain3 => mf20, bout0 => m19, bin0 => mf19, aout3 => m20, bin1 => mf18, aout2 => m21, bin2 => mf17, aout1 => m22, bin3 => mf16, aout0 => m23, benb => mfdrive);
  mf_1a23 : ic_74s241 port map(aenb_n => \-mfdrive\, ain0 => mf15, bout3 => m8, ain1 => mf14, bout2 => m9, ain2 => mf13, bout1 => m10, ain3 => mf12, bout0 => m11, bin0 => mf11, aout3 => m12, bin1 => mf10, aout2 => m13, bin2 => mf9, aout1 => m14, bin3 => mf8, aout0 => m15, benb => mfdrive);
  mf_1a25 : ic_74s241 port map(aenb_n => \-mfdrive\, ain0 => mf7, bout3 => m0, ain1 => mf6, bout2 => m1, ain2 => mf5, bout1 => m2, ain3 => mf4, bout0 => m3, bin0 => mf3, aout3 => m4, bin1 => mf2, aout2 => m5, bin2 => mf1, aout1 => m6, bin3 => mf0, aout0 => m7, benb => mfdrive);
  mf_1b24 : ic_74s241 port map(aenb_n => \-mfdrive\, ain0 => mf31, bout3 => m24, ain1 => mf30, bout2 => m25, ain2 => mf29, bout1 => m26, ain3 => mf28, bout0 => m27, bin0 => mf27, aout3 => m28, bin1 => mf26, aout2 => m29, bin2 => mf25, aout1 => m30, bin3 => mf24, aout0 => m31, benb => mfdrive);
  mf_2a04 : ic_74s08 port map(g2b     => tse1a, g2a => mfenb, g2q => mfdrive, g1b => '0', g1a => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  mf_3f14 : ic_74s02 port map(g3b     => pdlenb, g3a => spcenb, g3q_n => internal22, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4b => '0', g4a => '0');
  mf_4d06 : ic_74s08 port map(g4q     => mfenb, g4a => internal22, g4b => \-srcm\, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3a => '0', g3b => '0');
  mf_4d08 : ic_74s00 port map(g4q_n   => \-srcm\, g4a => \-ir31\, g4b=>\-mpass\, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0', g3b=>'0', g3a=>'0');

  --- Stack Buffer

  pdlptr_3c21 : ic_74s169 port map(up_dn  => \-srcpdlpop\, clk => clk3f, i0 => ob8, i1 => ob9, i2 => nc237, i3 => nc238, enb_p_n => gnd, load_n => \-destpdlp\, enb_t_n=>\-pdlcry7\, o3=>nc239, o2=>nc240, o1=>pdlptr9, o0=>pdlptr8, co_n=>nc241);
  pdlptr_3c22 : ic_25s07 port map(enb_n   => \-destpdlx\, d0 => pdlidx6, i0 => ob6, i1 => ob7, d1 => pdlidx7, i2 => ob8, d2 => pdlidx8, clk => clk3f, d3 => pdlidx9, i3 => ob9, d4 => nc233, i4 => nc234, i5 => nc235, d5 => nc236);
  pdlptr_3d24 : ic_74s169 port map(up_dn  => \-srcpdlpop\, clk => clk3f, i0 => ob4, i1 => ob5, i2 => ob6, i3 => ob7, enb_p_n => gnd, load_n => \-destpdlp\, enb_t_n=>\-pdlcry3\, o3=>pdlptr7, o2=>pdlptr6, o1=>pdlptr5, o0=>pdlptr4, co_n=>\-pdlcry7\);
  pdlptr_3d25 : ic_25s07 port map(enb_n   => \-destpdlx\, d0 => pdlidx0, i0 => ob0, i1 => ob1, d1 => pdlidx1, i2 => ob2, d2 => pdlidx2, clk => clk3f, d3 => pdlidx3, i3 => ob3, d4 => pdlidx4, i4 => ob4, i5 => ob5, d5 => pdlidx5);
  pdlptr_3d30 : ic_74s169 port map(up_dn  => \-srcpdlpop\, clk => clk3f, i0 => ob0, i1 => ob1, i2 => ob2, i3 => ob3, enb_p_n => gnd, load_n => \-destpdlp\, enb_t_n=>\-pdlcnt\, o3=>pdlptr3, o2=>pdlptr2, o1=>pdlptr1, o0=>pdlptr0, co_n=>\-pdlcry3\);
  pdlptr_4c01 : ic_74s241 port map(aenb_n => \-ppdrive\, ain0 => pdlptr3, bout3 => mf0, ain1 => pdlptr2, bout2 => mf1, ain2 => pdlptr1, bout1 => mf2, ain3 => pdlptr0, bout0 => mf3, bin0 => pdlidx3, aout3 => mf0, bin1 => pdlidx2, aout2 => mf1, bin2 => pdlidx1, aout1 => mf2, bin3 => pdlidx0, aout0 => mf3, benb => pidrive);
  pdlptr_4d04 : ic_74s241 port map(aenb_n => \-ppdrive\, ain0 => gnd, bout3 => mf8, ain1 => gnd, bout2 => mf9, ain2 => pdlptr9, bout1 => mf10, ain3 => pdlptr8, bout0 => mf11, bin0 => gnd, aout3 => mf8, bin1 => gnd, aout2 => mf9, bin2 => pdlidx9, aout1 => mf10, bin3 => pdlidx8, aout0 => mf11, benb => pidrive);
  pdlptr_4d05 : ic_74s241 port map(aenb_n => \-ppdrive\, ain0 => pdlptr7, bout3 => mf4, ain1 => pdlptr6, bout2 => mf5, ain2 => pdlptr5, bout1 => mf6, ain3 => pdlptr4, bout0 => mf7, bin0 => pdlidx7, aout3 => mf4, bin1 => pdlidx6, aout2 => mf5, bin2 => pdlidx5, aout1 => mf6, bin3 => pdlidx4, aout0 => mf7, benb => pidrive);
  pdlptr_4d06 : ic_74s08 port map(g3q     => pidrive, g3a => srcpdlidx, g3b => tse4b, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  pdlptr_4d08 : ic_74s00 port map(g3q_n   => \-ppdrive\, g3b => srcpdlptr, g3a => tse4b, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');

  pdlctl_4c11 : ic_74s175 port map(clr_n => \-reset\, q0 => pdlwrited, q0_n => \-pdlwrited\, d0=>pdlwrite, d1=>\-destpdl(x)\, q1_n=>pwidx, q1=>\-pwidx\, clk=>clk4f, q2=>imodd, q2_n=>\-imodd\, d2=>imod, d3=>\-destspc\, q3_n=>nc242, q3=>\-destspcd\);
  pdlctl_4c12 : ic_74s258 port map(sel   => \-pdlpb\, d0 => pdlptr0, d1 => pdlidx0, dy => \-pdla0b\, c0=>pdlptr1, c1=>pdlidx1, cy=>\-pdla1b\, by=>\-pdla2b\, b1=>pdlidx2, b0=>pdlptr2, ay=>\-pdla3b\, a1=>pdlidx3, a0=>pdlptr3, enb_n=>gnd);
  pdlctl_4c16 : ic_74s258 port map(sel   => \-pdlpa\, d0 => pdlptr8, d1 => pdlidx8, dy => \-pdla8b\, c0=>pdlptr9, c1=>pdlidx9, cy=>\-pdla9b\, by=>\-pdla0a\, b1=>pdlidx0, b0=>pdlptr0, ay=>\-pdla1a\, a1=>pdlidx1, a0=>pdlptr1, enb_n=>gnd);
  pdlctl_4c22 : ic_74s258 port map(sel   => \-pdlpa\, d0 => pdlptr2, d1 => pdlidx2, dy => \-pdla2a\, c0=>pdlptr3, c1=>pdlidx3, cy=>\-pdla3a\, by=>\-pdla4a\, b1=>pdlidx4, b0=>pdlptr4, ay=>\-pdla5a\, a1=>pdlidx5, a0=>pdlptr5, enb_n=>gnd);
  pdlctl_4d06 : ic_74s08 port map(g2b    => internal19, g2a => \-destpdl(p)\, g2q => \-pdlcnt\, g1b=>'0', g1a=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  pdlctl_4d07 : ic_74s51 port map(g1a    => \-pwidx\, g2a => clk4b, g2b => ir30, g2c => \-clk4e\, g2d=>\-pwidx\, g2y=>\-pdlpa\, g1y=>\-pdlpb\, g1c=>clk4b, g1d=>ir30, g1b=>\-clk4e\);
  pdlctl_4d08 : ic_74s00 port map(g1b    => \-srcpdlpop\, g1a => \-srcpdltop\, g1q_n=>pdlenb, g2b=>pdlenb, g2a=>tse4b, g2q_n=>\-pdldrive\, g3b=>'0', g3a=>'0', g4a=>'0', g4b=>'0');
  pdlctl_4d10 : ic_74s10 port map(g1a    => \-destpdltop\, g1b => \-destpdl(x)\, g1y_n=>pdlwrite, g1c=>\-destpdl(p)\, g2a=>'0', g2b=>'0', g2c=>'0', g3a=>'0', g3b=>'0', g3c=>'0');
  pdlctl_4d14 : ic_74s258 port map(sel   => \-pdlpb\, d0 => pdlptr4, d1 => pdlidx4, dy => \-pdla4b\, c0=>pdlptr5, c1=>pdlidx5, cy=>\-pdla5b\, by=>\-pdla6b\, b1=>pdlidx6, b0=>pdlptr6, ay=>\-pdla7b\, a1=>pdlidx7, a0=>pdlptr7, enb_n=>gnd);
  pdlctl_4d20 : ic_74s37 port map(g1a    => pdlwrited, g1b => wp4a, g1y => \-pwpa\, g2a => pdlwrited, g2b => wp4a, g2y => \-pwpb\, g3y=>\-pwpc\, g3a=>wp4a, g3b=>pdlwrited, g4a=>'0', g4b=>'0');
  pdlctl_4d24 : ic_74s258 port map(sel   => \-pdlpa\, d0 => pdlptr6, d1 => pdlidx6, dy => \-pdla6a\, c0=>pdlptr7, c1=>pdlidx7, cy=>\-pdla7a\, by=>\-pdla8a\, b1=>pdlidx8, b0=>pdlptr8, ay=>\-pdla9a\, a1=>pdlidx9, a0=>pdlptr9, enb_n=>gnd);
  pdlctl_4e03 : ic_74s32 port map(g3y    => internal19, g3a => \-srcpdlpop\, g3b => nop, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4a => '0', g4b => '0');

  pdl0_4c10 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdlparity, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>lparity);
  pdl0_4c13 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl28, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l28);
  pdl0_4c14 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl27, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l27);
  pdl0_4c15 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl26, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l26);
  pdl0_4c17 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl21, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpb\, di=>l21);
  pdl0_4c18 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl20, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpb\, di=>l20);
  pdl0_4c19 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl19, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpb\, di=>l19);
  pdl0_4c20 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl18, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpb\, di=>l18);
  pdl0_4d11 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl31, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l31);
  pdl0_4d12 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl30, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l30);
  pdl0_4d13 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl29, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l29);
  pdl0_4d16 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl25, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l25);
  pdl0_4d17 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl24, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l24);
  pdl0_4d18 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl23, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l23);
  pdl0_4d19 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl22, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpa\, di=>l22);
  pdl0_4d21 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl17, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpb\, di=>l17);
  pdl0_4d22 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0b\, a1 => \-pdla1b\, a2=>\-pdla2b\, a3=>\-pdla3b\, a4=>\-pdla4b\, do=>pdl16, a5=>\-pdla5b\, a6=>\-pdla6b\, a7=>\-pdla7b\, a8=>\-pdla8b\, a9=>\-pdla9b\, we_n=>\-pwpb\, di=>l16);

  pdl1_4c21 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl13, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpb\, di=>l13);
  pdl1_4c23 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl12, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpb\, di=>l12);
  pdl1_4c24 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl11, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpb\, di=>l11);
  pdl1_4c25 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl10, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l10);
  pdl1_4c26 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl4, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l4);
  pdl1_4c27 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl3, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l3);
  pdl1_4c28 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl2, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l2);
  pdl1_4c29 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl1, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l1);
  pdl1_4c30 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl0, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l0);
  pdl1_4d23 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl15, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpb\, di=>l15);
  pdl1_4d25 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl14, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpb\, di=>l14);
  pdl1_4d26 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl9, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l9);
  pdl1_4d27 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl8, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l8);
  pdl1_4d28 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl7, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l7);
  pdl1_4d29 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl6, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l6);
  pdl1_4d30 : ic_93425a port map(ce_n => gnd, a0 => \-pdla0a\, a1 => \-pdla1a\, a2=>\-pdla2a\, a3=>\-pdla3a\, a4=>\-pdla4a\, do=>pdl5, a5=>\-pdla5a\, a6=>\-pdla6a\, a7=>\-pdla7a\, a8=>\-pdla8a\, a9=>\-pdla9a\, we_n=>\-pwpc\, di=>l5);

  platch_4a02 : ic_74s373 port map(oenb_n => \-pdldrive\, o0 => m15, i0 => pdl15, i1 => pdl14, o1 => m14, o2 => m13, i2 => pdl13, i3 => pdl12, o3 => m12, hold_n => clk4a, o4 => m11, i4 => pdl11, i5 => pdl10, o5 => m10, o6 => m9, i6 => pdl9, i7 => pdl8, o7 => m8);
  platch_4a04 : ic_74s373 port map(oenb_n => \-pdldrive\, o0 => m7, i0 => pdl7, i1 => pdl6, o1 => m6, o2 => m5, i2 => pdl5, i3 => pdl4, o3 => m4, hold_n => clk4a, o4 => m3, i4 => pdl3, i5 => pdl2, o5 => m2, o6 => m1, i6 => pdl1, i7 => pdl0, o7 => m0);
  platch_4b03 : ic_74s373 port map(oenb_n => \-pdldrive\, o0 => m31, i0 => pdl31, i1 => pdl30, o1 => m30, o2 => m29, i2 => pdl29, i3 => pdl28, o3 => m28, hold_n => clk4a, o4 => m27, i4 => pdl27, i5 => pdl26, o5 => m26, o6 => m25, i6 => pdl25, i7 => pdl24, o7 => m24);
  platch_4b05 : ic_74s373 port map(oenb_n => \-pdldrive\, o0 => m23, i0 => pdl23, i1 => pdl22, o1 => m22, o2 => m21, i2 => pdl21, i3 => pdl20, o3 => m20, hold_n => clk4a, o4 => m19, i4 => pdl19, i5 => pdl18, o5 => m18, o6 => m17, i6 => pdl17, i7 => pdl16, o7 => m16);
  platch_4b08 : ic_74s373 port map(oenb_n => \-pdldrive\, o0 => nc219, i0 => nc220, i1 => nc221, o1 => nc222, o2 => nc223, i2 => nc224, i3 => nc225, o3 => nc226, hold_n => clk4a, o4 => nc227, i4 => nc228, i5 => nc229, o5 => nc230, o6 => nc231, i6 => nc232, i7 => pdlparity, o7 => mparity);

  --- The Shifter\Masker

  smctl_2d15 : ic_74s32 port map(g1a   => \-sh4\, g1b => \-sr\, g1y=>\-s4\, g2a=>'0', g2b=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  smctl_2d20 : ic_74s02 port map(g1q_n => \-mr\, g1a => \-irbyte\, g1b=>ir13, g2q_n=>\-sr\, g2a=>\-irbyte\, g2b=>ir12, g3b=>\-ir0\, g3a=>\-sr\, g3q_n=>s0, g4b=>\-ir1\, g4a=>\-sr\, g4q_n=>s1);
  smctl_2e10 : ic_74s283 port map(s1   => nc209, b1 => nc210, a1 => nc211, s0 => mskl4, a0 => ir9, b0 => mskr4, c0 => mskl3cry, c4 => nc212, s3 => nc213, b3 => nc214, a3 => nc215, s2 => nc216, a2 => nc217, b2 => nc218);
  smctl_2e14 : ic_74s02 port map(g1q_n => s3a, g1a => \-sr\, g1b => \-sh3\, g2q_n=>s3b, g2a=>\-sh3\, g2b=>\-sr\, g3b=>\-ir2\, g3a=>\-sr\, g3q_n=>s2a, g4b=>\-sr\, g4a=>\-ir2\, g4q_n=>s2b);
  smctl_2e19 : ic_74s02 port map(g1q_n => s4, g1a => \-sr\, g1b => \-sh4\, g2q_n=>mskr0, g2a=>\-mr\, g2b=>\-ir0\, g3b=>\-ir1\, g3a=>\-mr\, g3q_n=>mskr1, g4b=>\-ir2\, g4a=>\-mr\, g4q_n=>mskr2);
  smctl_2e25 : ic_74s283 port map(s1   => mskl1, b1 => mskr1, a1 => ir6, s0 => mskl0, a0 => ir5, b0 => mskr0, c0 => gnd, c4 => mskl3cry, s3 => mskl3, b3 => mskr3, a3 => ir8, s2 => mskl2, a2 => ir7, b2 => mskr2);
  smctl_2e30 : ic_74s02 port map(g1q_n => mskr3, g1a => \-mr\, g1b => \-sh3\, g2q_n=>mskr4, g2a=>\-mr\, g2b=>\-sh4\, g3b=>'0', g3a=>'0', g4b=>'0', g4a=>'0');

  shift0_2c21 : ic_25s10 port map(i_3 => m5, i_2 => m6, i_1 => m7, i0 => m8, i1 => m9, i2 => m10, i3 => m11, sel1 => s1, sel0 => s0, o3 => sa11, o2 => sa10, ce_n => gnd, o1 => sa9, o0 => sa8);
  shift0_2c26 : ic_25s10 port map(i_3 => m29, i_2 => m30, i_1 => m31, i0 => m0, i1 => m1, i2 => m2, i3 => m3, sel1 => s1, sel0 => s0, o3 => sa3, o2 => sa2, ce_n => gnd, o1 => sa1, o0 => sa0);
  shift0_2d25 : ic_25s10 port map(i_3 => m9, i_2 => m10, i_1 => m11, i0 => m12, i1 => m13, i2 => m14, i3 => m15, sel1 => s1, sel0 => s0, o3 => sa15, o2 => sa14, ce_n => gnd, o1 => sa13, o0 => sa12);
  shift0_2d30 : ic_25s10 port map(i_3 => m1, i_2 => m2, i_1 => m3, i0 => m4, i1 => m5, i2 => m6, i3 => m7, sel1 => s1, sel0 => s0, o3 => sa7, o2 => sa6, ce_n => gnd, o1 => sa5, o0 => sa4);
  shift0_2e21 : ic_25s10 port map(i_3 => sa6, i_2 => sa10, i_1 => sa14, i0 => sa18, i1 => sa22, i2 => sa26, i3 => sa30, sel1 => s3a, sel0 => s2a, o3 => r14, o2 => r10, ce_n => \-s4\, o1 => r6, o0 => r2);
  shift0_2e22 : ic_25s10 port map(i_3 => sa22, i_2 => sa26, i_1 => sa30, i0 => sa2, i1 => sa6, i2 => sa10, i3 => sa14, sel1 => s3a, sel0 => s2a, o3 => r14, o2 => r10, ce_n => s4, o1 => r6, o0 => r2);
  shift0_2e23 : ic_25s10 port map(i_3 => sa7, i_2 => sa11, i_1 => sa15, i0 => sa19, i1 => sa23, i2 => sa27, i3 => sa31, sel1 => s3a, sel0 => s2a, o3 => r15, o2 => r11, ce_n => \-s4\, o1 => r7, o0 => r3);
  shift0_2e24 : ic_25s10 port map(i_3 => sa23, i_2 => sa27, i_1 => sa31, i0 => sa3, i1 => sa7, i2 => sa11, i3 => sa15, sel1 => s3a, sel0 => s2a, o3 => r15, o2 => r11, ce_n => s4, o1 => r7, o0 => r3);
  shift0_2e26 : ic_25s10 port map(i_3 => sa4, i_2 => sa8, i_1 => sa12, i0 => sa16, i1 => sa20, i2 => sa24, i3 => sa28, sel1 => s3a, sel0 => s2a, o3 => r12, o2 => r8, ce_n => \-s4\, o1 => r4, o0 => r0);
  shift0_2e27 : ic_25s10 port map(i_3 => sa20, i_2 => sa24, i_1 => sa28, i0 => sa0, i1 => sa4, i2 => sa8, i3 => sa12, sel1 => s3a, sel0 => s2a, o3 => r12, o2 => r8, ce_n => s4, o1 => r4, o0 => r0);
  shift0_2e28 : ic_25s10 port map(i_3 => sa5, i_2 => sa9, i_1 => sa13, i0 => sa17, i1 => sa21, i2 => sa25, i3 => sa29, sel1 => s3a, sel0 => s2a, o3 => r13, o2 => r9, ce_n => \-s4\, o1 => r5, o0 => r1);
  shift0_2e29 : ic_25s10 port map(i_3 => sa21, i_2 => sa25, i_1 => sa29, i0 => sa1, i1 => sa5, i2 => sa9, i3 => sa13, sel1 => s3a, sel0 => s2a, o3 => r13, o2 => r9, ce_n => s4, o1 => r5, o0 => r1);

  shift1_2c01 : ic_25s10 port map(i_3 => m21, i_2 => m22, i_1 => m23, i0 => m24, i1 => m25, i2 => m26, i3 => m27, sel1 => s1, sel0 => s0, o3 => sa27, o2 => sa26, ce_n => gnd, o1 => sa25, o0 => sa24);
  shift1_2c06 : ic_25s10 port map(i_3 => m13, i_2 => m14, i_1 => m15, i0 => m16, i1 => m17, i2 => m18, i3 => m19, sel1 => s1, sel0 => s0, o3 => sa19, o2 => sa18, ce_n => gnd, o1 => sa17, o0 => sa16);
  shift1_2d05 : ic_25s10 port map(i_3 => m25, i_2 => m26, i_1 => m27, i0 => m28, i1 => m29, i2 => m30, i3 => m31, sel1 => s1, sel0 => s0, o3 => sa31, o2 => sa30, ce_n => gnd, o1 => sa29, o0 => sa28);
  shift1_2d10 : ic_25s10 port map(i_3 => m17, i_2 => m18, i_1 => m19, i0 => m20, i1 => m21, i2 => m22, i3 => m23, sel1 => s1, sel0 => s0, o3 => sa23, o2 => sa22, ce_n => gnd, o1 => sa21, o0 => sa20);
  shift1_2e01 : ic_25s10 port map(i_3 => sa22, i_2 => sa26, i_1 => sa30, i0 => sa2, i1 => sa6, i2 => sa10, i3 => sa14, sel1 => s3b, sel0 => s2b, o3 => r30, o2 => r26, ce_n => \-s4\, o1 => r22, o0 => r18);
  shift1_2e02 : ic_25s10 port map(i_3 => sa6, i_2 => sa10, i_1 => sa14, i0 => sa18, i1 => sa22, i2 => sa26, i3 => sa30, sel1 => s3b, sel0 => s2b, o3 => r30, o2 => r26, ce_n => s4, o1 => r22, o0 => r18);
  shift1_2e03 : ic_25s10 port map(i_3 => sa23, i_2 => sa27, i_1 => sa31, i0 => sa3, i1 => sa7, i2 => sa11, i3 => sa15, sel1 => s3b, sel0 => s2b, o3 => r31, o2 => r27, ce_n => \-s4\, o1 => r23, o0 => r19);
  shift1_2e04 : ic_25s10 port map(i_3 => sa7, i_2 => sa11, i_1 => sa15, i0 => sa19, i1 => sa23, i2 => sa27, i3 => sa31, sel1 => s3b, sel0 => s2b, o3 => r31, o2 => r27, ce_n => s4, o1 => r23, o0 => r19);
  shift1_2e06 : ic_25s10 port map(i_3 => sa20, i_2 => sa24, i_1 => sa28, i0 => sa0, i1 => sa4, i2 => sa8, i3 => sa12, sel1 => s3b, sel0 => s2b, o3 => r28, o2 => r24, ce_n => \-s4\, o1 => r20, o0 => r16);
  shift1_2e07 : ic_25s10 port map(i_3 => sa4, i_2 => sa8, i_1 => sa12, i0 => sa16, i1 => sa20, i2 => sa24, i3 => sa28, sel1 => s3b, sel0 => s2b, o3 => r28, o2 => r24, ce_n => s4, o1 => r20, o0 => r16);
  shift1_2e08 : ic_25s10 port map(i_3 => sa21, i_2 => sa25, i_1 => sa29, i0 => sa1, i1 => sa5, i2 => sa9, i3 => sa13, sel1 => s3b, sel0 => s2b, o3 => r29, o2 => r25, ce_n => \-s4\, o1 => r21, o0 => r17);
  shift1_2e09 : ic_25s10 port map(i_3 => sa5, i_2 => sa9, i_1 => sa13, i0 => sa17, i1 => sa21, i2 => sa25, i3 => sa29, sel1 => s3b, sel0 => s2b, o3 => r29, o2 => r25, ce_n => s4, o1 => r21, o0 => r17);

  mskg4_2d11 : ic_5600 port map(o0   => msk24, o1 => msk25, o2 => msk26, o3 => msk27, o4 => msk28, o5 => msk29, o6 => msk30, o7 => msk31, a0 => mskl0, a1 => mskl1, a2 => mskl2, a3 => mskl3, a4 => mskl4, ce_n => gnd);
  mskg4_2d12 : ic_5600 port map(o0   => msk24, o1 => msk25, o2 => msk26, o3 => msk27, o4 => msk28, o5 => msk29, o6 => msk30, o7 => msk31, a0 => mskr0, a1 => mskr1, a2 => mskr2, a3 => mskr3, a4 => mskr4, ce_n => gnd);
  mskg4_2d16 : ic_5600 port map(o0   => msk8, o1 => msk9, o2 => msk10, o3 => msk11, o4 => msk12, o5 => msk13, o6 => msk14, o7 => msk15, a0 => mskl0, a1 => mskl1, a2 => mskl2, a3 => mskl3, a4 => mskl4, ce_n => gnd);
  mskg4_2d17 : ic_5600 port map(o0   => msk8, o1 => msk9, o2 => msk10, o3 => msk11, o4 => msk12, o5 => msk13, o6 => msk14, o7 => msk15, a0 => mskr0, a1 => mskr1, a2 => mskr2, a3 => mskr3, a4 => mskr4, ce_n => gnd);
  mskg4_2d26 : ic_74s04 port map(g1a => nc253, g1q_n => nc254, g2a => ir31, g2q_n => \-ir31\, g3a => ir13, g3q_n => \-ir13\, g4q=>\-ir12\, g4a=>ir12, g5q_n=>nc255, g5a=>nc256, g6q_n=>nc257, g6a=>nc258);
  mskg4_2e11 : ic_5600 port map(o0   => msk16, o1 => msk17, o2 => msk18, o3 => msk19, o4 => msk20, o5 => msk21, o6 => msk22, o7 => msk23, a0 => mskl0, a1 => mskl1, a2 => mskl2, a3 => mskl3, a4 => mskl4, ce_n => gnd);
  mskg4_2e12 : ic_5600 port map(o0   => msk16, o1 => msk17, o2 => msk18, o3 => msk19, o4 => msk20, o5 => msk21, o6 => msk22, o7 => msk23, a0 => mskr0, a1 => mskr1, a2 => mskr2, a3 => mskr3, a4 => mskr4, ce_n => gnd);
  mskg4_2e15 : ic_res20 port map(r2  => aeqm, r3 => msk31, r4 => msk30, r5 => msk29, r6 => msk28, r7 => msk27, r8 => msk26, r9 => msk25, r11 => msk24, r12 => msk23, r13 => msk22, r14 => msk21, r15 => msk20, r16 => msk19, r17 => msk18, r18 => msk17, r19 => msk16, r10 => '0');
  mskg4_2e16 : ic_5600 port map(o0   => msk0, o1 => msk1, o2 => msk2, o3 => msk3, o4 => msk4, o5 => msk5, o6 => msk6, o7 => msk7, a0 => mskl0, a1 => mskl1, a2 => mskl2, a3 => mskl3, a4 => mskl4, ce_n => gnd);
  mskg4_2e17 : ic_5600 port map(o0   => msk0, o1 => msk1, o2 => msk2, o3 => msk3, o4 => msk4, o5 => msk5, o6 => msk6, o7 => msk7, a0 => mskr0, a1 => mskr1, a2 => mskr2, a3 => mskr3, a4 => mskr4, ce_n => gnd);
  mskg4_2e20 : ic_res20 port map(r2  => nc252, r3 => msk15, r4 => msk14, r5 => msk13, r6 => msk12, r7 => msk11, r8 => msk10, r9 => msk9, r11 => msk8, r12 => msk7, r13 => msk6, r14 => msk5, r15 => msk4, r16 => msk3, r17 => msk2, r18 => msk1, r19 => msk0, r10 => '0');

  --- The ALU

  aluc4_2a16 : ic_74s37 port map(g1a     => \-aluf0\, g1b => \-aluf0\, g1y=>aluf0b, g2a=>\-aluf1\, g2b=>\-aluf1\, g2y=>aluf1b, g3y=>aluf2b, g3a=>\-aluf2\, g3b=>\-aluf2\, g4y=>aluf3b, g4a=>\-aluf3\, g4b=>\-aluf3\);
  aluc4_2a17 : ic_74s37 port map(g1a     => \-aluf0\, g1b => \-aluf0\, g1y=>aluf0a, g2a=>\-aluf1\, g2b=>\-aluf1\, g2y=>aluf1a, g3y=>aluf2a, g3a=>\-aluf2\, g3b=>\-aluf2\, g4y=>aluf3a, g4a=>\-aluf3\, g4b=>\-aluf3\);
  aluc4_2a18 : ic_74s182 port map(y1     => yy1, x1 => xx1, y0 => yy0, x0 => xx0, y3 => nc437, x3 => nc438, xout => nc439, cout2_n => nc440, yout => nc441, cout1_n => \-cin32\, cout0_n => \-cin16\, cin_n=>\-cin0\, y2=>nc442, x2=>nc443);
  aluc4_2a19 : ic_74s182 port map(y1     => yout23, x1 => xout23, y0 => yout19, x0 => xout19, y3 => yout31, x3 => xout31, xout => xx1, cout2_n => \-cin28\, yout => yy1, cout1_n => \-cin24\, cout0_n=>\-cin20\, cin_n=>\-cin16\, y2=>yout27, x2=>xout27);
  aluc4_2a20 : ic_74s182 port map(y1     => yout7, x1 => xout7, y0 => yout3, x0 => xout3, y3 => yout15, x3 => xout15, xout => xx0, cout2_n => \-cin12\, yout => yy0, cout1_n => \-cin8\, cout0_n=>\-cin4\, cin_n=>\-cin0\, y2=>yout11, x2=>xout11);
  aluc4_2b16 : ic_74s153 port map(enb1_n => gnd, sel1 => alusub, g1c3 => gnd, g1c2 => hi12, g1c1 => gnd, g1c0 => \-ir3\, g1q => \-aluf3\, g2q=>\-aluf2\, g2c0=>\-ir4\, g2c1=>hi12, g2c2=>gnd, g2c3=>gnd, sel0=>aluadd, enb2_n=>gnd);
  aluc4_2b17 : ic_74s153 port map(enb1_n => gnd, sel1 => alusub, g1c3 => gnd, g1c2 => gnd, g1c1 => hi12, g1c0 => ir6, g1q => \-aluf1\, g2q => \-aluf0\, g2c0=>ir5, g2c1=>gnd, g2c2=>hi12, g2c3=>gnd, sel0=>aluadd, enb2_n=>gnd);
  aluc4_2b18 : ic_74s153 port map(enb1_n => gnd, sel1 => alusub, g1c3 => gnd, g1c2 => hi12, g1c1 => hi12, g1c0 => ir7, g1q => \-alumode\, g2q => \-cin0\, g2c0=>\-ir2\, g2c1=>hi12, g2c2=>irjump, g2c3=>gnd, sel0=>aluadd, enb2_n=>gnd);
  aluc4_2b20 : ic_74s37 port map(g1a     => \-alumode\, g1b => \-alumode\, g1y=>alumode, g2a=>'0', g2b=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  aluc4_2c10 : ic_74s02 port map(g1q_n   => internal33, g1a => ir5, g1b => \-divposlasttime\, g2q_n => \-divposlasttime\, g2a=>q0, g2b=>ir6, g3b=>\-divposlasttime\, g3a=>\-div\, g3q_n=>divsubcond, g4b=>internal33, g4a=>\-div\, g4q_n=>divaddcond);
  aluc4_2c11 : ic_74s04 port map(g1a     => a31b, g1q_n => \-a31\, g2a => ir4, g2q_n => \-ir4\, g3a=>ir3, g3q_n=>\-ir3\, g4q=>\-ir2\, g4a=>ir2, g5q_n=>\-ir1\, g5a=>ir1, g6q_n=>\-ir0\, g6a=>ir0);
  aluc4_2c15 : ic_74s00 port map(g1b     => divaddcond, g1a => \-a31\, g1q_n => internal34, g2b => divsubcond, g2a => a31a, g2q_n => internal35, g3q_n => internal36, g3b => divsubcond, g3a => \-a31\, g4q_n=>internal37, g4a=>divaddcond, g4b=>a31a);
  aluc4_2c20 : ic_74s20 port map(g1a     => \-mulnop\, g1b => internal36, g1c => internal37, g1d => \-irjump\, g1y_n=>alusub, g2y_n=>aluadd, g2a=>\-mul\, g2b=>hi12, g2c=>internal35, g2d=>internal34);
  aluc4_2d15 : ic_74s32 port map(g2a     => \-mul\, g2b => q0, g2y => \-mulnop\, g1a=>'0', g1b=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  aluc4_2d21 : ic_7428 port map(g1q_n    => osel1a, g1a => \-ir13\, g1b => \-iralu\, g2q_n=>osel0a, g2a=>\-ir12\, g2b=>\-iralu\, g3a=>\-iralu\, g3b=>\-ir13\, g3q_n=>osel1b, g4a=>\-iralu\, g4b=>\-ir12\, g4q_n=>osel0b);

  alu0_2a23 : ic_74s181 port map(b0 => a12, a0 => m12, s3 => aluf3b, s2 => aluf2b, s1 => aluf1b, s0 => aluf0b, cin_n => \-cin12\, m => alumode, f0 => alu12, f1 => alu13, f2 => alu14, f3 => alu15, aeb => aeqm, x => xout15, cout_n => nc461, y => yout15, b3 => a15, a3 => m15, b2 => a14, a2 => m14, b1 => a13, a1 => m13);
  alu0_2a28 : ic_74s181 port map(b0 => a4, a0 => m4, s3 => aluf3b, s2 => aluf2b, s1 => aluf1b, s0 => aluf0b, cin_n => \-cin4\, m => alumode, f0 => alu4, f1 => alu5, f2 => alu6, f3 => alu7, aeb => aeqm, x => xout7, cout_n => nc463, y => yout7, b3 => a7, a3 => m7, b2 => a6, a2 => m6, b1 => a5, a1 => m5);
  alu0_2b23 : ic_74s181 port map(b0 => a8, a0 => m8, s3 => aluf3b, s2 => aluf2b, s1 => aluf1b, s0 => aluf0b, cin_n => \-cin8\, m => alumode, f0 => alu8, f1 => alu9, f2 => alu10, f3 => alu11, aeb => aeqm, x => xout11, cout_n => nc462, y => yout11, b3 => a11, a3 => m11, b2 => a10, a2 => m10, b1 => a9, a1 => m9);
  alu0_2b28 : ic_74s181 port map(b0 => a0, a0 => m0, s3 => aluf3b, s2 => aluf2b, s1 => aluf1b, s0 => aluf0b, cin_n => \-cin0\, m => alumode, f0 => alu0, f1 => alu1, f2 => alu2, f3 => alu3, aeb => aeqm, x => xout3, cout_n => nc464, y => yout3, b3 => a3, a3 => m3, b2 => a2, a2 => m2, b1 => a1, a1 => m1);

  alu1_2a03 : ic_74s181 port map(b0 => a31a, a0 => m31b, s3 => aluf3a, s2 => aluf2a, s1 => aluf1a, s0 => aluf0a, cin_n => \-cin32\, m => alumode, f0 => alu32, f1 => nc444, f2 => nc445, f3 => nc446, aeb => nc447, x => nc448, cout_n => nc449, y => nc450, b3 => nc451, a3 => nc452, b2 => nc453, a2 => nc454, b1 => nc455, a1 => nc456);
  alu1_2a04 : ic_74s08 port map(g1b => m31, g1a => hi12, g1q => m31b, g2b => '0', g2a => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  alu1_2a08 : ic_74s181 port map(b0 => a28, a0 => m28, s3 => aluf3a, s2 => aluf2a, s1 => aluf1a, s0 => aluf0a, cin_n => \-cin28\, m => alumode, f0 => alu28, f1 => alu29, f2 => alu30, f3 => alu31, aeb => aeqm, x => xout31, cout_n => nc457, y => yout31, b3 => a31b, a3 => m31b, b2 => a30, a2 => m30, b1 => a29, a1 => m29);
  alu1_2a13 : ic_74s181 port map(b0 => a20, a0 => m20, s3 => aluf3a, s2 => aluf2a, s1 => aluf1a, s0 => aluf0a, cin_n => \-cin20\, m => alumode, f0 => alu20, f1 => alu21, f2 => alu22, f3 => alu23, aeb => aeqm, x => xout23, cout_n => nc459, y => yout23, b3 => a23, a3 => m23, b2 => a22, a2 => m22, b1 => a21, a1 => m21);
  alu1_2b08 : ic_74s181 port map(b0 => a24, a0 => m24, s3 => aluf3a, s2 => aluf2a, s1 => aluf1a, s0 => aluf0a, cin_n => \-cin24\, m => alumode, f0 => alu24, f1 => alu25, f2 => alu26, f3 => alu27, aeb => aeqm, x => xout27, cout_n => nc458, y => yout27, b3 => a27, a3 => m27, b2 => a26, a2 => m26, b1 => a25, a1 => m25);
  alu1_2b13 : ic_74s181 port map(b0 => a16, a0 => m16, s3 => aluf3a, s2 => aluf2a, s1 => aluf1a, s0 => aluf0a, cin_n => \-cin16\, m => alumode, f0 => alu16, f1 => alu17, f2 => alu18, f3 => alu19, aeb => aeqm, x => xout19, cout_n => nc460, y => yout19, b3 => a19, a3 => m19, b2 => a18, a2 => m18, b1 => a17, a1 => m17);

  --- The Q Register

  qctl_1a18 : ic_74s00 port map(g3q_n   => \-qdrive\, g3b => tse2, g3a => srcq, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  qctl_1e12 : ic_74s241 port map(aenb_n => \-qdrive\, ain0 => q7, bout3 => mf0, ain1 => q6, bout2 => mf1, ain2 => q5, bout1 => mf2, ain3 => q4, bout0 => mf3, bin0 => q3, aout3 => mf4, bin1 => q2, aout2 => mf5, bin2 => q1, aout1 => mf6, bin3 => q0, aout0 => mf7, benb => qdrive);
  qctl_1f08 : ic_74s241 port map(aenb_n => \-qdrive\, ain0 => q31, bout3 => mf24, ain1 => q30, bout2 => mf25, ain2 => q29, bout1 => mf26, ain3 => q28, bout0 => mf27, bin0 => q27, aout3 => mf28, bin1 => q26, aout2 => mf29, bin2 => q25, aout1 => mf30, bin3 => q24, aout0 => mf31, benb => qdrive);
  qctl_1f10 : ic_74s241 port map(aenb_n => \-qdrive\, ain0 => q23, bout3 => mf16, ain1 => q22, bout2 => mf17, ain2 => q21, bout1 => mf18, ain3 => q20, bout0 => mf19, bin0 => q19, aout3 => mf20, bin1 => q18, aout2 => mf21, bin2 => q17, aout1 => mf22, bin3 => q16, aout0 => mf23, benb => qdrive);
  qctl_1f15 : ic_74s241 port map(aenb_n => \-qdrive\, ain0 => q15, bout3 => mf8, ain1 => q14, bout2 => mf9, ain2 => q13, bout1 => mf10, ain3 => q12, bout0 => mf11, bin0 => q11, aout3 => mf12, bin1 => q10, aout2 => mf13, bin2 => q9, aout1 => mf14, bin3 => q8, aout0 => mf15, benb => qdrive);
  qctl_2a04 : ic_74s08 port map(g4q     => qdrive, g4a => tse2, g4b => srcq, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3a => '0', g3b => '0');
  qctl_2a05 : ic_74s04 port map(g5q_n   => srcq, g5a => \-srcq\, g6q_n => \-alu31\, g6a=>alu31, g1a=>'0', g2a=>'0', g3a=>'0', g4a=>'0');
  qctl_2b19 : ic_7428 port map(g3a      => \-iralu\, g3b => \-ir1\, g3q_n=>qs1, g4a=>\-iralu\, g4b=>\-ir0\, g4q_n=>qs0, g1a=>'0', g1b=>'0', g2a=>'0', g2b=>'0');

  q_2c07 : ic_74s194 port map(clr_n => hi7, sir => q23, i0 => alu24, i1 => alu25, i2 => alu26, i3 => alu27, sil => q28, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q27, q2 => q26, q1 => q25, q0 => q24);
  q_2c08 : ic_74s194 port map(clr_n => hi7, sir => q27, i0 => alu28, i1 => alu29, i2 => alu30, i3 => alu31, sil => alu0, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q31, q2 => q30, q1 => q29, q0 => q28);
  q_2c12 : ic_74s194 port map(clr_n => hi7, sir => q15, i0 => alu16, i1 => alu17, i2 => alu18, i3 => alu19, sil => q20, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q19, q2 => q18, q1 => q17, q0 => q16);
  q_2c13 : ic_74s194 port map(clr_n => hi7, sir => q19, i0 => alu20, i1 => alu21, i2 => alu22, i3 => alu23, sil => q24, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q23, q2 => q22, q1 => q21, q0 => q20);
  q_2c22 : ic_74s194 port map(clr_n => hi7, sir => q7, i0 => alu8, i1 => alu9, i2 => alu10, i3 => alu11, sil => q12, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q11, q2 => q10, q1 => q9, q0 => q8);
  q_2c23 : ic_74s194 port map(clr_n => hi7, sir => q11, i0 => alu12, i1 => alu13, i2 => alu14, i3 => alu15, sil => q16, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q15, q2 => q14, q1 => q13, q0 => q12);
  q_2c27 : ic_74s194 port map(clr_n => hi7, sir => \-alu31\, i0 => alu0, i1 => alu1, i2 => alu2, i3 => alu3, sil => q4, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q3, q2 => q2, q1 => q1, q0 => q0);
  q_2c28 : ic_74s194 port map(clr_n => hi7, sir => q3, i0 => alu4, i1 => alu5, i2 => alu6, i3 => alu7, sil => q8, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q7, q2 => q6, q1 => q5, q0 => q4);

  --- The L Register

  l_3c26 : ic_74s374 port map(oenb_n => gnd, o0 => l7, i0 => ob7, i1 => ob6, o1 => l6, o2 => l5, i2 => ob5, i3 => ob4, o3 => l4, clk => clk3f, o4 => l3, i4 => ob3, i5 => ob2, o5 => l2, o6 => l1, i6 => ob1, i7 => ob0, o7 => l0);
  l_3c27 : ic_74s374 port map(oenb_n => gnd, o0 => l15, i0 => ob15, i1 => ob14, o1 => l14, o2 => l13, i2 => ob13, i3 => ob12, o3 => l12, clk => clk3f, o4 => l11, i4 => ob11, i5 => ob10, o5 => l10, o6 => l9, i6 => ob9, i7 => ob8, o7 => l8);
  l_3c28 : ic_74s374 port map(oenb_n => gnd, o0 => l23, i0 => ob23, i1 => ob22, o1 => l22, o2 => l21, i2 => ob21, i3 => ob20, o3 => l20, clk => clk3f, o4 => l19, i4 => ob19, i5 => ob18, o5 => l18, o6 => l17, i6 => ob17, i7 => ob16, o7 => l16);
  l_3c29 : ic_74s374 port map(oenb_n => gnd, o0 => l31, i0 => ob31, i1 => ob30, o1 => l30, o2 => l29, i2 => ob29, i3 => ob28, o3 => l28, clk => clk3f, o4 => l27, i4 => ob27, i5 => ob26, o5 => l26, o6 => l25, i6 => ob25, i7 => ob24, o7 => l24);
  l_4c03 : ic_93s48 port map(i6      => l5, i5 => l6, i4 => l7, i3 => l8, i2 => l9, i1 => l10, i0 => l11, po => lparl, pe => nc369, i11 => l0, i10 => l1, i9 => l2, i8 => l3, i7 => l4);
  l_4c08 : ic_93s48 port map(i6      => l17, i5 => l18, i4 => l19, i3 => l20, i2 => l21, i1 => l22, i0 => l23, po => nc370, pe => \-lparm\, i11 => l12, i10 => l13, i9 => l14, i8 => l15, i7 => l16);
  l_4c09 : ic_93s48 port map(i6      => l25, i5 => l26, i4 => l27, i3 => l28, i2 => l29, i1 => l30, i0 => l31, po => lparity, pe => \-lparity\, i11 => lparl, i10 => \-lparm\, i9=>gnd, i8=>gnd, i7=>l24);

  --- The Dispatch Memory

  dspctl_2f22 : ic_5610 port map(o0       => dmask0, o1 => dmask1, o2 => dmask2, o3 => dmask3, o4 => dmask4, o5 => dmask5, o6 => dmask6, o7 => nc407, a0 => ir5, a1 => ir6, a2 => ir7, a3 => gnd, a4 => gnd, ce_n => gnd);
  dspctl_3c14 : ic_25s07 port map(enb_n   => \-irdisp\, d0 => dc6, i0 => ir38, i1 => ir39, d1 => dc7, i2 => ir40, d2 => dc8, clk => clk3e, d3 => dc9, i3 => ir41, d4 => nc403, i4 => nc404, i5 => nc405, d5 => nc406);
  dspctl_3c15 : ic_25s07 port map(enb_n   => \-irdisp\, d0 => dc0, i0 => ir32, i1 => ir33, d1 => dc1, i2 => ir34, d2 => dc2, clk => clk3e, d3 => dc3, i3 => ir35, d4 => dc4, i4 => ir36, i5 => ir37, d5 => dc5);
  dspctl_3d02 : ic_74s00 port map(g1b     => dpareven, g1a => dispenb, g1q_n => dparok, g2b => '0', g2a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  dspctl_3e19 : ic_74s86 port map(g3y     => dpareven, g3a => \-dparh\, g3b => dparl, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4a => '0', g4b => '0');
  dspctl_3f11 : ic_74s241 port map(aenb_n => hi4, ain0 => nc389, bout3 => aa16, ain1 => nc390, bout2 => aa17, ain2 => nc391, bout1 => nc392, ain3 => nc393, bout0 => nc394, bin0 => nc395, aout3 => nc396, bin1 => nc397, aout2 => nc398, bin2 => a17, aout1 => nc399, bin3 => a16, aout0 => nc400, benb => hi4);
  dspctl_3f12 : ic_74s241 port map(aenb_n => gnd, ain0 => a15, bout3 => aa8, ain1 => a14, bout2 => aa9, ain2 => a13, bout1 => aa10, ain3 => a12, bout0 => aa11, bin0 => a11, aout3 => aa12, bin1 => a10, aout2 => aa13, bin2 => a9, aout1 => aa14, bin3 => a8, aout0 => aa15, benb => hi4);
  dspctl_3f13 : ic_74s241 port map(aenb_n => gnd, ain0 => a7, bout3 => aa0, ain1 => a6, bout2 => aa1, ain2 => a5, bout1 => aa2, ain3 => a4, bout0 => aa3, bin0 => a3, aout3 => aa4, bin1 => a2, aout2 => aa5, bin2 => a1, aout1 => aa6, bin3 => a0, aout0 => aa7, benb => hi4);
  dspctl_3f14 : ic_74s02 port map(g1q_n   => \-dmapbenb\, g1a => ir8, g1b => ir9, g2q_n => dispwr, g2a => \-irdisp\, g2b=>\-funct2\, g3b=>'0', g3a=>'0', g4b=>'0', g4a=>'0');
  dspctl_4f09 : ic_74s280 port map(i0     => dpc9, i1 => dpc10, i2 => dpc11, even => \-dparh\, odd => nc402, i3 => dpc12, i4 => dpc13, i5 => dn, i6 => dp, i7 => dr, i8 => dpar);
  dspctl_4f10 : ic_74s280 port map(i0     => dpc0, i1 => dpc1, i2 => dpc2, even => nc401, odd => dparl, i3 => dpc3, i4 => dpc4, i5 => dpc5, i6 => dpc6, i7 => dpc7, i8 => dpc8);

  dram0_2f03 : ic_74s37 port map(g1a     => wp2, g1b => dispwr, g1y => \-dwea\, g2a => '0', g2b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  dram0_2f21 : ic_74s04 port map(g1a     => nc418, g1q_n => nc419, g2a => \-dadr10a\, g2q_n => dadr10a, g3a => ir22b, g3q_n => \-dadr10a\, g4q=>\-dadr9a\, g4a=>ir21b, g5q_n=>\-dadr8a\, g5a=>ir20b, g6q_n=>\-dadr7a\, g6a=>ir19b);
  dram0_2f24 : ic_74s64 port map(d4      => ir12b, b2 => vmo19, a2 => ir9b, c3 => r0, b3 => dmask0, a3 => \-dmapbenb\, \out\=>\-dadr0a\, a1 => vmo18, b1 => ir8b, c4 => hi6, b4 => hi6, a4 => hi6);
  dram0_2f25 : ic_74s241 port map(aenb_n => gnd, ain0 => ir12, bout3 => ir19b, ain1 => ir13, bout2 => ir18b, ain2 => ir14, bout1 => ir17b, ain3 => ir15, bout0 => ir16b, bin0 => ir16, aout3 => ir15b, bin1 => ir17, aout2 => ir14b, bin2 => ir18, aout1 => ir13b, bin3 => ir19, aout0 => ir12b, benb => hi6);
  dram0_2f26 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc5, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa5);
  dram0_2f27 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1=>\-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc5, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa5);
  dram0_2f28 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc4, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa4);
  dram0_2f29 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1=>\-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc4, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa4);
  dram0_2f30 : ic_74s51 port map(g1a     => r3, g2a => ir18b, g2b => hi6, g2c => dmask6, g2d => r6, g2y => \-dadr6a\, g1y => \-dadr3a\, g1c=>ir15b, g1d=>hi6, g1b=>dmask3);
  dram0_3f01 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc3, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa3);
  dram0_3f02 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1=>\-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc3, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa3);
  dram0_3f03 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc2, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa2);
  dram0_3f04 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1=>\-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc2, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa2);
  dram0_3f05 : ic_74s51 port map(g1a     => r2, g2a => ir17b, g2b => hi4, g2c => dmask5, g2d => r5, g2y => \-dadr5a\, g1y => \-dadr2a\, g1c=>ir14b, g1d=>hi4, g1b=>dmask2);
  dram0_3f06 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc1, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa1);
  dram0_3f07 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1=>\-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc1, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa1);
  dram0_3f08 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0a\, a1 => \-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc0, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa0);
  dram0_3f09 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0a\, a1=>\-dadr1a\, a2=>\-dadr2a\, a3=>\-dadr3a\, a4=>\-dadr4a\, do=>dpc0, a5=>\-dadr5a\, a6=>\-dadr6a\, a7=>\-dadr7a\, a8=>\-dadr8a\, a9=>\-dadr9a\, we_n=>\-dwea\, di=>aa0);
  dram0_3f10 : ic_74s51 port map(g1a     => r1, g2a => ir16b, g2b => hi4, g2c => dmask4, g2d => r4, g2y => \-dadr4a\, g1y => \-dadr1a\, g1c=>ir13b, g1d=>hi4, g1b=>dmask1);

  dram1_2f03 : ic_74s37 port map(g2a     => wp2, g2b => dispwr, g2y => \-dweb\, g1a => '0', g1b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  dram1_2f04 : ic_74s04 port map(g1a     => nc416, g1q_n => nc417, g2a => \-vmo19\, g2q_n => vmo19, g3a => \-vmo18\, g3q_n=>vmo18, g4q=>\-dadr9b\, g4a=>ir21b, g5q_n=>\-dadr8b\, g5a=>ir20b, g6q_n=>\-dadr7b\, g6a=>ir19b);
  dram1_2f05 : ic_74s64 port map(d4      => ir12b, b2 => vmo19, a2 => ir9b, c3 => r0, b3 => dmask0, a3 => \-dmapbenb\, \out\=>\-dadr0b\, a1 => vmo18, b1 => ir8b, c4 => hi6, b4 => hi6, a4 => hi6);
  dram1_2f06 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0b\, a1 => \-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc11, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa11);
  dram1_2f07 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0b\, a1=>\-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc11, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa11);
  dram1_2f08 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0b\, a1 => \-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc10, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa10);
  dram1_2f09 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0b\, a1=>\-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc10, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa10);
  dram1_2f10 : ic_74s51 port map(g1a     => r3, g2a => ir18b, g2b => hi6, g2c => dmask6, g2d => r6, g2y => \-dadr6b\, g1y => \-dadr3b\, g1c=>ir15b, g1d=>hi6, g1b=>dmask3);
  dram1_2f11 : ic_93425a port map(ce_n   => dadr10a, a0 => \-dadr0b\, a1 => \-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc9, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa9);
  dram1_2f12 : ic_93425a port map(ce_n   => \-dadr10a\, a0 => \-dadr0b\, a1=>\-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc9, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa9);
  dram1_2f13 : ic_93425a port map(ce_n   => dadr10c, a0 => \-dadr0b\, a1 => \-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc8, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa8);
  dram1_2f14 : ic_93425a port map(ce_n   => \-dadr10c\, a0 => \-dadr0b\, a1=>\-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc8, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa8);
  dram1_2f15 : ic_74s51 port map(g1a     => r2, g2a => ir17b, g2b => hi6, g2c => dmask5, g2d => r5, g2y => \-dadr5b\, g1y => \-dadr2b\, g1c=>ir14b, g1d=>hi6, g1b=>dmask2);
  dram1_2f16 : ic_93425a port map(ce_n   => dadr10c, a0 => \-dadr0b\, a1 => \-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc7, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa7);
  dram1_2f17 : ic_93425a port map(ce_n   => \-dadr10c\, a0 => \-dadr0b\, a1=>\-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc7, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa7);
  dram1_2f18 : ic_93425a port map(ce_n   => dadr10c, a0 => \-dadr0b\, a1 => \-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc6, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa6);
  dram1_2f19 : ic_93425a port map(ce_n   => \-dadr10c\, a0 => \-dadr0b\, a1=>\-dadr1b\, a2=>\-dadr2b\, a3=>\-dadr3b\, a4=>\-dadr4b\, do=>dpc6, a5=>\-dadr5b\, a6=>\-dadr6b\, a7=>\-dadr7b\, a8=>\-dadr8b\, a9=>\-dadr9b\, we_n=>\-dweb\, di=>aa6);
  dram1_2f20 : ic_74s51 port map(g1a     => r1, g2a => ir16b, g2b => hi6, g2c => dmask4, g2d => r4, g2y => \-dadr4b\, g1y => \-dadr1b\, g1c=>ir13b, g1d=>hi6, g1b=>dmask1);
  dram1_2f23 : ic_74s241 port map(aenb_n => gnd, ain0 => ir20, bout3 => nc410, ain1 => ir21, bout2 => nc411, ain2 => ir22, bout1 => nc412, ain3 => ir8, bout0 => ir9b, bin0 => ir9, aout3 => ir8b, bin1 => nc413, aout2 => ir22b, bin2 => nc414, aout1 => ir21b, bin3 => nc415, aout0 => ir20b, benb => hi6);

  dram2_1f16 : ic_93425a port map(ce_n => dadr10c, a0 => \-dadr0c\, a1 => \-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dpar, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa17);
  dram2_1f17 : ic_93425a port map(ce_n => \-dadr10c\, a0 => \-dadr0c\, a1=>\-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dpar, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa17);
  dram2_1f18 : ic_93425a port map(ce_n => dadr10c, a0 => \-dadr0c\, a1 => \-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dr, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa16);
  dram2_1f19 : ic_93425a port map(ce_n => \-dadr10c\, a0 => \-dadr0c\, a1=>\-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dr, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa16);
  dram2_1f20 : ic_74s51 port map(g1a   => r3, g2a => ir18b, g2b => hi11, g2c => dmask6, g2d => r6, g2y => \-dadr6c\, g1y => \-dadr3c\, g1c=>ir15b, g1d=>hi11, g1b=>dmask3);
  dram2_1f21 : ic_93425a port map(ce_n => dadr10c, a0 => \-dadr0c\, a1 => \-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dp, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa15);
  dram2_1f22 : ic_93425a port map(ce_n => \-dadr10c\, a0 => \-dadr0c\, a1=>\-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dp, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa15);
  dram2_1f23 : ic_93425a port map(ce_n => dadr10c, a0 => \-dadr0c\, a1 => \-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dn, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa14);
  dram2_1f24 : ic_93425a port map(ce_n => \-dadr10c\, a0 => \-dadr0c\, a1=>\-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dn, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa14);
  dram2_1f25 : ic_74s51 port map(g1a   => r2, g2a => ir17b, g2b => hi11, g2c => dmask5, g2d => r5, g2y => \-dadr5c\, g1y => \-dadr2c\, g1c=>ir14b, g1d=>hi11, g1b=>dmask2);
  dram2_1f26 : ic_93425a port map(ce_n => dadr10c, a0 => \-dadr0c\, a1 => \-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dpc13, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa13);
  dram2_1f27 : ic_93425a port map(ce_n => \-dadr10c\, a0 => \-dadr0c\, a1=>\-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dpc13, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa13);
  dram2_1f28 : ic_93425a port map(ce_n => dadr10c, a0 => \-dadr0c\, a1 => \-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dpc12, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa12);
  dram2_1f29 : ic_93425a port map(ce_n => \-dadr10c\, a0 => \-dadr0c\, a1=>\-dadr1c\, a2=>\-dadr2c\, a3=>\-dadr3c\, a4=>\-dadr4c\, do=>dpc12, a5=>\-dadr5c\, a6=>\-dadr6c\, a7=>\-dadr7c\, a8=>\-dadr8c\, a9=>\-dadr9c\, we_n=>\-dwec\, di=>aa12);
  dram2_1f30 : ic_74s51 port map(g1a   => r1, g2a => ir16b, g2b => hi11, g2c => dmask4, g2d => r4, g2y => \-dadr4c\, g1y => \-dadr1c\, g1c=>ir13b, g1d=>hi11, g1b=>dmask1);
  dram2_2f01 : ic_74s64 port map(d4    => ir12b, b2 => vmo19, a2 => ir9b, c3 => r0, b3 => dmask0, a3 => \-dmapbenb\, \out\=>\-dadr0c\, a1 => vmo18, b1 => ir8b, c4 => hi6, b4 => hi6, a4 => hi6);
  dram2_2f02 : ic_74s04 port map(g1a   => nc408, g1q_n => nc409, g2a => \-dadr10c\, g2q_n => dadr10c, g3a => ir22b, g3q_n => \-dadr10c\, g4q=>\-dadr9c\, g4a=>ir21b, g5q_n=>\-dadr8c\, g5a=>ir20b, g6q_n=>\-dadr7c\, g6a=>ir19b);
  dram2_2f03 : ic_74s37 port map(g3y   => \-dwec\, g3a => dispwr, g3b => wp2, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4a => '0', g4b => '0');

  --- Jump Conditions

  flag_3e07 : ic_74s00 port map(g1b   => ir45, g1a => \-nopa\, g1q_n => \-ilong\, g2b=>'0', g2a=>'0', g3b=>'0', g3a=>'0', g4a=>'0', g4b=>'0');
  flag_3e08 : ic_25ls2519 port map(i0 => ob29, q0a => nc385, q0b => \lc_byte_mode\, i1 => ob28, q1a => nc386, q1b => \prog.unibus.reset\, o_enb_n=>hi4, out_enb_n=>gnd, clk=>clk3c, q2b=>\int.enable\, q2a=>nc387, i2=>ob27, q3b=>\sequence.break\, q3a=>nc388, i3=>ob26, clk_enb_n=>\-destintctl\, inv=>hi4, asyn_clr_n=>\-reset\);
  flag_3e11 : ic_74s00 port map(g4q_n => \-statbit\, g4a => \-nopa\, g4b=>ir46, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0', g3b=>'0', g3a=>'0');
  flag_3e13 : ic_74s151 port map(i3   => aeqm, i2 => alu32, i1 => aluneg, i0 => r0, q => jcond, q_n => \-jcond\, ce_n => gnd, sel2 => conds2, sel1 => conds1, sel0 => conds0, i7 => hi4, i6 => \pgf.or.int.or.sb\, i5=>\pgf.or.int\, i4=>\-vmaok\);
  flag_3e14 : ic_74s08 port map(g1b   => ir2, g1a => ir5, g1q => conds2, g2b => ir1, g2a => ir5, g2q => conds1, g3q => conds0, g3a => ir5, g3b => ir0, g4a => '0', g4b => '0');
  flag_3e17 : ic_74s02 port map(g4b   => \-alu32\, g4a => aeqm, g4q_n => aluneg, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g3b => '0', g3a => '0');
  flag_3e18 : ic_74s32 port map(g2a   => \-vmaok\, g2b => sint, g2y => \pgf.or.int\, g3y=>internal30, g3a=>\sequence.break\, g3b=>sint, g4y=>\pgf.or.int.or.sb\, g4a=>internal30, g4b=>\-vmaok\, g1a=>'0', g1b=>'0');
  flag_3e22 : ic_74s04 port map(g4q   => \-alu32\, g4a => alu32, g1a => '0', g2a => '0', g3a => '0', g5a => '0', g6a => '0');
  flag_4d09 : ic_74s08 port map(g3q   => sint, g3a => \int.enable\, g3b => sintr, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');

  --- Flow of Control

  contrl_3d21 : ic_74s08 port map(g1b    => spushd, g1a => tse3a, g1q => spcwpass, g2b => \-ipopj\, g2a => \-iwrited\, g2q=>\-popj\, g3q=>spcdrive, g3a=>spcenb, g3b=>tse3a, g4a=>'0', g4b=>'0');
  contrl_3d26 : ic_74s175 port map(clr_n => \-reset\, q0 => inop, q0_n => \-inop\, d0=>n, d1=>nc420, q1_n=>nc421, q1=>nc422, clk=>clk3c, q2=>spushd, q2_n=>\-spushd\, d2=>spush, d3=>iwrite, q3_n=>\-iwrited\, q3=>iwrited);
  contrl_3d28 : ic_74s00 port map(g1b    => \-srcspc\, g1a => \-srcspcpop\, g1q_n=>spcenb, g2b=>spcenb, g2a=>tse3a, g2q_n=>\-spcdrive\, g3q_n=>\-spcpass\, g3b=>tse3a, g3a=>\-spushd\, g4q_n=>\-spcwpass\, g4a=>tse3a, g4b=>spushd);
  contrl_3e07 : ic_74s00 port map(g2b    => ir42, g2a => \-nop\, g2q_n => \-ipopj\, g1b=>'0', g1a=>'0', g3b=>'0', g3a=>'0', g4a=>'0', g4b=>'0');
  contrl_3e09 : ic_74s32 port map(g1a    => \-srcspcpop\, g1b => nop, g1y => \-srcspcpopreal\, g2a=>'0', g2b=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  contrl_3e14 : ic_74s08 port map(g4q    => \-nopa\, g4a => \-nop11\, g4b=>\-inop\, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0', g3a=>'0', g3b=>'0');
  contrl_3e18 : ic_74s32 port map(g1a    => \-irdisp\, g1b => dr, g1y => \-ignpopj\, g2a=>'0', g2b=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  contrl_3e22 : ic_74s04 port map(g1a    => \-destspc\, g1q_n => destspc, g2a => nop, g2q_n => \-nop\, g3a=>'0', g4a=>'0', g5a=>'0', g6a=>'0');
  contrl_3e23 : ic_74s00 port map(g1b    => dr, g1a => dp, g1q_n => \-dfall\, g2b => \-trap\, g2a=>internal32, g2q_n=>n, g3q_n=>internal31, g3b=>\-popj\, g3a=>\-srcspcpopreal\, g4q_n=>nop, g4a=>\-trap\, g4b=>\-nopa\);
  contrl_3e24 : ic_74s08 port map(g1b    => irdisp, g1a => \-funct2\, g1q => dispenb, g2b => irjump, g2a => ir6, g2q => jfalse, g3q => jcalf, g3a => ir8, g3b => jfalse, g4q => jretf, g4a => ir6, g4b => jret);
  contrl_3e25 : ic_74s64 port map(d4     => ir7, b2 => dn, a2 => dispenb, c3 => ir7, b3 => \-jcond\, a3 => jfalse, \out\=>internal32, a1 => hi4, b1 => iwrited, c4 => jcond, b4 => \-ir6\, a4=>irjump);
  contrl_3e26 : ic_74s64 port map(d4     => jcond, b2 => \-jcond\, a2 => jcalf, c3 => \-dr\, b3=>dp, a3=>dispenb, \out\=>\-spush\, a1=>hi4, b1=>destspc, c4=>ir8, b4=>\-ir6\, a4=>irjump);
  contrl_3e27 : ic_74s64 port map(d4     => hi4, b2 => \-jcond\, a2 => jfalse, c3 => jcond, b3 => \-ir6\, a3=>irjump, \out\=>pcs1, a1=>\-ignpopj\, b1=>popj, c4=>\-dp\, b4=>dr, a4=>dispenb);
  contrl_3e28 : ic_74s64 port map(d4     => hi4, b2 => \-jcond\, a2 => jretf, c3 => jcond, b3 => \-ir6\, a3=>jret, \out\=>\-spop\, a1=>\-ignpopj\, b1=>internal31, c4=>\-dp\, b4=>dr, a4=>dispenb);
  contrl_3e29 : ic_74s11 port map(g1a    => \-ir8\, g1b => irjump, g2a => irjump, g2b => ir8, g2c => ir9, g2y_n => iwrite, g1y_n => jret, g1c => ir9, g3a => '0', g3b => '0', g3c => '0');
  contrl_3f20 : ic_74s04 port map(g1a    => \-popj\, g1q_n => popj, g2a => ir8, g2q_n => \-ir8\, g3a=>ir6, g3q_n=>\-ir6\, g4q=>spush, g4a=>\-spush\, g5q_n=>\-dp\, g5a=>dp, g6q_n=>\-dr\, g6a=>dr);
  contrl_3f30 : ic_74s64 port map(d4     => hi4, b2 => \-dfall\, a2 => dispenb, c3 => hi4, b3 => \-jcond\, a3=>jretf, \out\=>pcs0, a1=>hi4, b1=>popj, c4=>jcond, b4=>\-ir6\, a4=>jret);
  contrl_4d09 : ic_74s08 port map(g1b    => \-spush\, g1a => \-spop\, g1q=>\-spcnt\, g2b=>'0', g2a=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  contrl_4e30 : ic_74s37 port map(g1a    => \-destspcd\, g1b => \-destspcd\, g1y=>destspcd, g2a=>wp4c, g2b=>spushd, g2y=>\-swpb\, g3y=>\-swpa\, g3a=>spushd, g3b=>wp4c, g4a=>'0', g4b=>'0');

  --- Microcode Subroutine Return Stack

  spc_4e21 : ic_82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw14, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco14, d1 => spco15, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw15, we1_n => gnd);
  spc_4e22 : ic_82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw12, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco12, d1 => spco13, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw13, we1_n => gnd);
  spc_4e23 : ic_82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw10, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco10, d1 => spco11, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw11, we1_n => gnd);
  spc_4e24 : ic_res20 port map(r2     => spcopar, r3 => spco18, r4 => spco17, r5 => spco16, r6 => spco15, r7 => hi1, r8 => hi2, r9 => hi3, r11 => hi4, r12 => hi5, r13 => hi6, r14 => hi7, r15 => spco14, r16 => spco13, r17 => spco12, r18 => spco11, r19 => spco10, r10 => '0');
  spc_4e26 : ic_82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw4, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco4, d1 => spco5, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw5, we1_n => gnd);
  spc_4e27 : ic_82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw2, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco2, d1 => spco3, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw3, we1_n => gnd);
  spc_4e28 : ic_82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw0, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco0, d1 => spco1, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw1, we1_n => gnd);
  spc_4e29 : ic_res20 port map(r2     => spco9, r3 => spco8, r4 => spco7, r5 => spco6, r6 => spco5, r7 => hi8, r8 => hi9, r9 => hi10, r11 => hi11, r12 => hi12, r13 => nc182, r14 => nc183, r15 => spco4, r16 => spco3, r17 => spco2, r18 => spco1, r19 => spco0, r10 => '0');
  spc_4f23 : ic_74s169 port map(up_dn => spush, clk => clk4f, i0 => nc192, i1 => nc193, i2 => nc194, i3 => nc195, enb_p_n => gnd, load_n => hi1, enb_t_n => \-spcnt\, o3 => spcptr3, o2 => spcptr2, o1 => spcptr1, o0 => spcptr0, co_n => \-spccry\);
  spc_4f24 : ic_82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw18, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco18, d1 => spcopar, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcwpar, we1_n => gnd);
  spc_4f25 : ic_82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw16, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco16, d1 => spco17, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw17, we1_n => gnd);
  spc_4f28 : ic_74s169 port map(up_dn => spush, clk => clk4f, i0 => nc184, i1 => nc185, i2 => nc186, i3 => nc187, enb_p_n => gnd, load_n => hi1, enb_t_n => \-spccry\, o3 => nc188, o2 => nc189, o1 => nc190, o0 => spcptr4, co_n => nc191);
  spc_4f29 : ic_82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw8, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco8, d1 => spco9, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw9, we1_n => gnd);
  spc_4f30 : ic_82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw6, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco6, d1 => spco7, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw7, we1_n => gnd);

  spclch_4a07 : ic_74s373 port map(oenb_n => \-spcdrive\, o0 => m23, i0 => gnd, i1 => gnd, o1 => m22, o2 => m21, i2 => gnd, i3 => gnd, o3 => m20, hold_n => clk4c, o4 => m19, i4 => gnd, i5 => spco18, o5 => m18, o6 => m17, i6 => spco17, i7 => spco16, o7 => m16);
  spclch_4a09 : ic_74s373 port map(oenb_n => \-spcdrive\, o0 => m15, i0 => spco15, i1 => spco14, o1 => m14, o2 => m13, i2 => spco13, i3 => spco12, o3 => m12, hold_n => clk4c, o4 => m11, i4 => spco11, i5 => spco10, o5 => m10, o6 => m9, i6 => spco9, i7 => spco8, o7 => m8);
  spclch_4a10 : ic_74s373 port map(oenb_n => \-spcdrive\, o0 => m7, i0 => spco7, i1 => spco6, o1 => m6, o2 => m5, i2 => spco5, i3 => spco4, o3 => m4, hold_n => clk4c, o4 => m3, i4 => spco3, i5 => spco2, o5 => m2, o6 => m1, i6 => spco1, i7 => spco0, o7 => m0);
  spclch_4b10 : ic_74s241 port map(aenb_n => \-spcdrive\, ain0 => gnd, bout3 => m24, ain1 => gnd, bout2 => m25, ain2 => gnd, bout1 => m26, ain3 => spcptr4, bout0 => m27, bin0 => spcptr3, aout3 => m28, bin1 => spcptr2, aout2 => m29, bin2 => spcptr1, aout1 => m30, bin3 => spcptr0, aout0 => m31, benb => spcdrive);
  spclch_4e16 : ic_74s241 port map(aenb_n => hi1, ain0 => nc166, bout3 => spc16, ain1 => nc167, bout2 => spc17, ain2 => nc168, bout1 => spc18, ain3 => nc169, bout0 => spcpar, bin0 => spcwpar, aout3 => nc170, bin1 => spcw18, aout2 => nc171, bin2 => spcw17, aout1 => nc172, bin3 => spcw16, aout0 => nc173, benb => spcwpass);
  spclch_4e17 : ic_74s241 port map(aenb_n => \-spcwpass\, ain0 => spcw15, bout3 => spc8, ain1 => spcw14, bout2 => spc9, ain2 => spcw13, bout1 => spc10, ain3 => spcw12, bout0 => spc11, bin0 => spcw11, aout3 => spc12, bin1 => spcw10, aout2 => spc13, bin2 => spcw9, aout1 => spc14, bin3 => spcw8, aout0 => spc15, benb => spcwpass);
  spclch_4e18 : ic_74s241 port map(aenb_n => \-spcwpass\, ain0 => spcw7, bout3 => spc0, ain1 => spcw6, bout2 => spc1, ain2 => spcw5, bout1 => spc2, ain3 => spcw4, bout0 => spc3, bin0 => spcw3, aout3 => spc4, bin1 => spcw2, aout2 => spc5, bin2 => spcw1, aout1 => spc6, bin3 => spcw0, aout0 => spc7, benb => spcwpass);
  spclch_4f18 : ic_74s373 port map(oenb_n => \-spcpass\, o0 => nc174, i0 => nc175, i1 => nc176, o1 => nc177, o2 => nc178, i2 => nc179, i3 => nc180, o3 => nc181, hold_n => clk4d, o4 => spcpar, i4 => spcopar, i5 => spco18, o5 => spc18, o6 => spc17, i6 => spco17, i7 => spco16, o7 => spc16);
  spclch_4f19 : ic_74s373 port map(oenb_n => \-spcpass\, o0 => spc15, i0 => spco15, i1 => spco14, o1 => spc14, o2 => spc13, i2 => spco13, i3 => spco12, o3 => spc12, hold_n => clk4d, o4 => spc11, i4 => spco11, i5 => spco10, o5 => spc10, o6 => spc9, i6 => spco9, i7 => spco8, o7 => spc8);
  spclch_4f20 : ic_74s373 port map(oenb_n => \-spcpass\, o0 => spc7, i0 => spco7, i1 => spco6, o1 => spc6, o2 => spc5, i2 => spco5, i3 => spco4, o3 => spc4, hold_n => clk4d, o4 => spc3, i4 => spco3, i5 => spco2, o5 => spc2, o6 => spc1, i6 => spco1, i7 => spco0, o7 => spc0);

  spcw_4e11 : ic_74s157 port map(sel => destspcd, a4 => reta12, b4 => l12, y4 => spcw12, a3 => reta13, b3 => l13, y3 => spcw13, y2 => spcw14, b2 => l14, a2 => gnd, y1 => spcw15, b1 => l15, a1 => gnd, enb_n => gnd);
  spcw_4e12 : ic_74s157 port map(sel => destspcd, a4 => reta8, b4 => l8, y4 => spcw8, a3 => reta9, b3 => l9, y3 => spcw9, y2 => spcw10, b2 => l10, a2 => reta10, y1 => spcw11, b1 => l11, a1 => reta11, enb_n => gnd);
  spcw_4e13 : ic_74s157 port map(sel => destspcd, a4 => reta4, b4 => l4, y4 => spcw4, a3 => reta5, b3 => l5, y3 => spcw5, y2 => spcw6, b2 => l6, a2 => reta6, y1 => spcw7, b1 => l7, a1 => reta7, enb_n => gnd);
  spcw_4e14 : ic_74s157 port map(sel => destspcd, a4 => reta0, b4 => l0, y4 => spcw0, a3 => reta1, b3 => l1, y3 => spcw1, y2 => spcw2, b2 => l2, a2 => reta2, y1 => spcw3, b1 => l3, a1 => reta3, enb_n => gnd);
  spcw_4f11 : ic_25s09 port map(sel  => n, aq => reta12, a0 => ipc12, a1 => wpc12, b1 => wpc13, b0 => ipc13, bq => reta13, clk => clk4d, cq => nc153, c0 => nc154, c1 => nc155, d1 => nc156, d0 => nc157, dq => nc158);
  spcw_4f12 : ic_25s09 port map(sel  => n, aq => reta8, a0 => ipc8, a1 => wpc8, b1 => wpc9, b0 => ipc9, bq => reta9, clk => clk4d, cq => reta10, c0 => ipc10, c1 => wpc10, d1 => wpc11, d0 => ipc11, dq => reta11);
  spcw_4f13 : ic_25s09 port map(sel  => n, aq => reta4, a0 => ipc4, a1 => wpc4, b1 => wpc5, b0 => ipc5, bq => reta5, clk => clk4d, cq => reta6, c0 => ipc6, c1 => wpc6, d1 => wpc7, d0 => ipc7, dq => reta7);
  spcw_4f14 : ic_25s09 port map(sel  => n, aq => reta0, a0 => ipc0, a1 => wpc0, b1 => wpc1, b0 => ipc1, bq => reta1, clk => clk4d, cq => reta2, c0 => ipc2, c1 => wpc2, d1 => wpc3, d0 => ipc3, dq => reta3);
  spcw_4f15 : ic_74s157 port map(sel => destspcd, a4 => gnd, b4 => l16, y4 => spcw16, a3 => gnd, b3 => l17, y3 => spcw17, y2 => spcw18, b2 => l18, a2 => gnd, y1 => nc159, b1 => nc160, a1 => nc161, enb_n => gnd);

  spcpar_3e19 : ic_74s86 port map(g2a => spcwparh, g2b => \-spcwparl\, g2y => spcwpar, g1a => '0', g1b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  spcpar_4f16 : ic_93s48 port map(i6  => spcw17, i5 => spcw18, i4 => gnd, i3 => gnd, i2 => gnd, i1 => gnd, i0 => gnd, po => spcwparh, pe => nc162, i11 => spcw12, i10 => spcw13, i9 => spcw14, i8 => spcw15, i7 => spcw16);
  spcpar_4f17 : ic_93s48 port map(i6  => spcw5, i5 => spcw6, i4 => spcw7, i3 => spcw8, i2 => spcw9, i1 => spcw10, i0 => spcw11, po => nc163, pe => \-spcwparl\, i11 => spcw0, i10 => spcw1, i9 => spcw2, i8 => spcw3, i7 => spcw4);
  spcpar_4f21 : ic_93s48 port map(i6  => spc16, i5 => spc17, i4 => spc18, i3 => spcpar, i2 => gnd, i1 => gnd, i0 => gnd, po => spcparh, pe => nc164, i11 => spc11, i10 => spc12, i9 => spc13, i8 => spc14, i7 => spc15);
  spcpar_4f26 : ic_93s48 port map(i6  => spc5, i5 => spc6, i4 => spc7, i3 => spc8, i2 => spc9, i1 => spc10, i0 => spcparh, po => spcparok, pe => nc165, i11 => spc0, i10 => spc1, i9 => spc2, i8 => spc3, i7 => spc4);

  lpc_4d01 : ic_74s241 port map(aenb_n => gnd, ain0 => pc8, bout3 => nc341, ain1 => pc9, bout2 => nc342, ain2 => pc10, bout1 => pc13b, ain3 => pc11, bout0 => pc12b, bin0 => pc12, aout3 => pc11b, bin1 => pc13, aout2 => pc10b, bin2 => nc343, aout1 => pc9b, bin3 => nc344, aout0 => pc8b, benb => hi5);
  lpc_4d02 : ic_74s241 port map(aenb_n => gnd, ain0 => pc0, bout3 => pc7b, ain1 => pc1, bout2 => pc6b, ain2 => pc2, bout1 => pc5b, ain3 => pc3, bout0 => pc4b, bin0 => pc4, aout3 => pc3b, bin1 => pc5, aout2 => pc2b, bin2 => pc6, aout1 => pc1b, bin3 => pc7, aout0 => pc0b, benb => hi5);
  lpc_4d06 : ic_74s08 port map(g1b     => irdisp, g1a => ir25, g1q => internal23, g2b => '0', g2a => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  lpc_4e06 : ic_74s157 port map(sel    => internal23, a4 => pc12, b4 => lpc12, y4 => wpc12, a3 => pc13, b3 => lpc13, y3 => wpc13, y2 => nc345, b2 => nc346, a2 => nc347, y1 => nc348, b1 => nc349, a1 => nc350, enb_n => gnd);
  lpc_4e07 : ic_74s157 port map(sel    => internal24, a4 => pc8, b4 => lpc8, y4 => wpc8, a3 => pc9, b3 => lpc9, y3 => wpc9, y2 => wpc10, b2 => lpc10, a2 => pc10, y1 => wpc11, b1 => lpc11, a1 => pc11, enb_n => gnd);
  lpc_4e08 : ic_74s157 port map(sel    => internal24, a4 => pc4, b4 => lpc4, y4 => wpc4, a3 => pc5, b3 => lpc5, y3 => wpc5, y2 => wpc6, b2 => lpc6, a2 => pc6, y1 => wpc7, b1 => lpc7, a1 => pc7, enb_n => gnd);
  lpc_4e09 : ic_74s157 port map(sel    => internal24, a4 => pc0, b4 => lpc0, y4 => wpc0, a3 => pc1, b3 => lpc1, y3 => wpc1, y2 => wpc2, b2 => lpc2, a2 => pc2, y1 => wpc3, b1 => lpc3, a1 => pc3, enb_n => gnd);
  lpc_4f06 : ic_25s07 port map(enb_n   => \lpc.hold\, d0 => lpc5, i0 => pc5, i1 => pc4, d1 => lpc4, i2 => pc3, d2 => lpc3, clk => clk4b, d3 => lpc2, i3 => pc2, d4 => lpc1, i4 => pc1, i5 => pc0, d5 => lpc0);
  lpc_4f07 : ic_25s07 port map(enb_n   => \lpc.hold\, d0 => lpc11, i0 => pc11, i1 => pc10, d1 => lpc10, i2 => pc9, d2 => lpc9, clk => clk4b, d3 => lpc8, i3 => pc8, d4 => lpc7, i4 => pc7, i5 => pc6, d5 => lpc6);
  lpc_4f08 : ic_25s07 port map(enb_n   => \lpc.hold\, d0 => nc351, i0 => nc352, i1 => nc353, d1 => nc354, i2 => nc355, d2 => nc356, clk => clk4b, d3 => nc357, i3 => nc358, d4 => lpc13, i4 => pc13, i5 => pc12, d5 => lpc12);

  --- Next PC Selector

  npc_3f26 : ic_74s283 port map(s1     => ipc13, b1 => gnd, a1 => pc13, s0 => ipc12, a0 => pc12, b0 => gnd, c0 => pccry11, c4 => nc243, s3 => nc244, b3 => gnd, a3 => nc245, s2 => nc246, a2 => nc247, b2 => gnd);
  npc_3f27 : ic_74s283 port map(s1     => ipc9, b1 => gnd, a1 => pc9, s0 => ipc8, a0 => pc8, b0 => gnd, c0 => pccry7, c4 => pccry11, s3 => ipc11, b3 => gnd, a3 => pc11, s2 => ipc10, a2 => pc10, b2 => gnd);
  npc_3f28 : ic_74s283 port map(s1     => ipc5, b1 => gnd, a1 => pc5, s0 => ipc4, a0 => pc4, b0 => gnd, c0 => pccry3, c4 => pccry7, s3 => ipc7, b3 => gnd, a3 => pc7, s2 => ipc6, a2 => pc6, b2 => gnd);
  npc_3f29 : ic_74s283 port map(s1     => ipc1, b1 => gnd, a1 => pc1, s0 => ipc0, a0 => pc0, b0 => gnd, c0 => hi4, c4 => pccry3, s3 => ipc3, b3 => gnd, a3 => pc3, s2 => ipc2, a2 => pc2, b2 => gnd);
  npc_4e01 : ic_74s153 port map(enb1_n => trapb, sel1 => pcs1, g1c3 => ipc3, g1c2 => dpc3, g1c1 => ir15, g1c0 => spc3, g1q => npc3, g2q => npc2, g2c0 => spc2, g2c1 => ir14, g2c2 => dpc2, g2c3 => ipc2, sel0 => pcs0, enb2_n => trapb);
  npc_4e02 : ic_74s153 port map(enb1_n => trapb, sel1 => pcs1, g1c3 => ipc1, g1c2 => dpc1, g1c1 => ir13, g1c0 => spc1a, g1q => npc1, g2q => npc0, g2c0 => spc0, g2c1 => ir12, g2c2 => dpc0, g2c3 => ipc0, sel0 => pcs0, enb2_n => trapb);
  npc_4e04 : ic_74s374 port map(oenb_n => gnd, o0 => nc248, i0 => nc249, i1 => nc250, o1 => nc251, o2 => pc13, i2 => npc13, i3 => npc12, o3 => pc12, clk => clk4b, o4 => pc11, i4 => npc11, i5 => npc10, o5 => pc10, o6 => pc9, i6 => npc9, i7 => npc8, o7 => pc8);
  npc_4e05 : ic_74s374 port map(oenb_n => gnd, o0 => pc7, i0 => npc7, i1 => npc6, o1 => pc6, o2 => pc5, i2 => npc5, i3 => npc4, o3 => pc4, clk => clk4b, o4 => pc3, i4 => npc3, i5 => npc2, o5 => pc2, o6 => pc1, i6 => npc1, i7 => npc0, o7 => pc0);
  npc_4f01 : ic_74s153 port map(enb1_n => trapa, sel1 => pcs1, g1c3 => ipc13, g1c2 => dpc13, g1c1 => ir25, g1c0 => spc13, g1q => npc13, g2q => npc12, g2c0 => spc12, g2c1 => ir24, g2c2 => dpc12, g2c3 => ipc12, sel0 => pcs0, enb2_n => trapa);
  npc_4f02 : ic_74s153 port map(enb1_n => trapa, sel1 => pcs1, g1c3 => ipc11, g1c2 => dpc11, g1c1 => ir23, g1c0 => spc11, g1q => npc11, g2q => npc10, g2c0 => spc10, g2c1 => ir22, g2c2 => dpc10, g2c3 => ipc10, sel0 => pcs0, enb2_n => trapa);
  npc_4f03 : ic_74s153 port map(enb1_n => trapa, sel1 => pcs1, g1c3 => ipc9, g1c2 => dpc9, g1c1 => ir21, g1c0 => spc9, g1q => npc9, g2q => npc8, g2c0 => spc8, g2c1 => ir20, g2c2 => dpc8, g2c3 => ipc8, sel0 => pcs0, enb2_n => trapa);
  npc_4f04 : ic_74s153 port map(enb1_n => trapa, sel1 => pcs1, g1c3 => ipc7, g1c2 => dpc7, g1c1 => ir19, g1c0 => spc7, g1q => npc7, g2q => npc6, g2c0 => spc6, g2c1 => ir18, g2c2 => dpc6, g2c3 => ipc6, sel0 => pcs0, enb2_n => trapb);
  npc_4f05 : ic_74s153 port map(enb1_n => trapb, sel1 => pcs1, g1c3 => ipc5, g1c2 => dpc5, g1c1 => ir17, g1c0 => spc5, g1q => npc5, g2q => npc4, g2c0 => spc4, g2c1 => ir16, g2c2 => dpc4, g2c3 => ipc4, sel0 => pcs0, enb2_n => trapb);

  --- The LC register and Instruction Prefetch

  lc_1a16 : ic_74s241 port map(aenb_n => \-lcdrive\, ain0 => needfetch, bout3 => mf24, ain1 => gnd, bout2 => mf25, ain2 => \lc_byte_mode\, bout1=>mf26, ain3=>\prog.unibus.reset\, bout0=>mf27, bin0=>\int.enable\, aout3=>mf28, bin1=>\sequence.break\, aout2=>mf29, bin2=>lc25, aout1=>mf30, bin3=>lc24, aout0=>mf31, benb=>lcdrive);
  lc_1a18 : ic_74s00 port map(g2b     => srclc, g2a => tse1a, g2q_n => \-lcdrive\, g1b => '0', g1a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  lc_1a20 : ic_74s241 port map(aenb_n => \-lcdrive\, ain0 => lc7, bout3 => mf0, ain1 => lc6, bout2 => mf1, ain2 => lc5, bout1 => mf2, ain3 => lc4, bout0 => mf3, bin0 => lc3, aout3 => mf4, bin1 => lc2, aout2 => mf5, bin2 => lc1, aout1 => mf6, bin3 => lc0b, aout0 => mf7, benb => lcdrive);
  lc_1a22 : ic_74s241 port map(aenb_n => \-lcdrive\, ain0 => lc23, bout3 => mf16, ain1 => lc22, bout2 => mf17, ain2 => lc21, bout1 => mf18, ain3 => lc20, bout0 => mf19, bin0 => lc19, aout3 => mf20, bin1 => lc18, aout2 => mf21, bin2 => lc17, aout1 => mf22, bin3 => lc16, aout0 => mf23, benb => lcdrive);
  lc_1a24 : ic_74s241 port map(aenb_n => \-lcdrive\, ain0 => lc15, bout3 => mf8, ain1 => lc14, bout2 => mf9, ain2 => lc13, bout1 => mf10, ain3 => lc12, bout0 => mf11, bin0 => lc11, aout3 => mf12, bin1 => lc10, aout2 => mf13, bin2 => lc9, aout1 => mf14, bin3 => lc8, aout0 => mf15, benb => lcdrive);
  lc_1a26 : ic_74s169 port map(up_dn  => hi11, clk => clk1a, i0 => ob20, i1 => ob21, i2 => ob22, i3 => ob23, enb_p_n => gnd, load_n => \-destlc\, enb_t_n => \-lcry19\, o3=>lc23, o2=>lc22, o1=>lc21, o0=>lc20, co_n=>\-lcry23\);
  lc_1b28 : ic_74s169 port map(up_dn  => hi11, clk => clk1a, i0 => ob16, i1 => ob17, i2 => ob18, i3 => ob19, enb_p_n => gnd, load_n => \-destlc\, enb_t_n => \-lcry15\, o3=>lc19, o2=>lc18, o1=>lc17, o0=>lc16, co_n=>\-lcry19\);
  lc_1c30 : ic_74s169 port map(up_dn  => hi11, clk => clk2a, i0 => ob12, i1 => ob13, i2 => ob14, i3 => ob15, enb_p_n => gnd, load_n => \-destlc\, enb_t_n => \-lcry11\, o3=>lc15, o2=>lc14, o1=>lc13, o0=>lc12, co_n=>\-lcry15\);
  lc_1d29 : ic_74s169 port map(up_dn  => hi11, clk => clk2c, i0 => ob8, i1 => ob9, i2 => ob10, i3 => ob11, enb_p_n => gnd, load_n => \-destlc\, enb_t_n => \-lcry7\, o3=>lc11, o2=>lc10, o1=>lc9, o0=>lc8, co_n=>\-lcry11\);
  lc_2a04 : ic_74s08 port map(g3q     => lcdrive, g3a => tse1a, g3b => srclc, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  lc_2a05 : ic_74s04 port map(g1a     => \-srclc\, g1q_n => srclc, g2a => '0', g3a => '0', g4a => '0', g5a => '0', g6a => '0');
  lc_2b03 : ic_74s169 port map(up_dn  => hi11, clk => clk1a, i0 => ob24, i1 => ob25, i2 => nc364, i3 => nc365, enb_p_n => gnd, load_n => \-destlc\, enb_t_n => \-lcry23\, o3=>nc366, o2=>nc367, o1=>lc25, o0=>lc24, co_n=>nc368);
  lc_2c05 : ic_74s169 port map(up_dn  => hi11, clk => clk2a, i0 => ob4, i1 => ob5, i2 => ob6, i3 => ob7, enb_p_n => gnd, load_n => \-destlc\, enb_t_n => \-lcry3\, o3=>lc7, o2=>lc6, o1=>lc5, o0=>lc4, co_n=>\-lcry7\);

  lcc_1c15 : ic_74s02 port map(g3b    => \lc_byte_mode\, g3a => \-lcinc\, g3q_n=>internal25, g1a=>'0', g1b=>'0', g2a=>'0', g2b=>'0', g4b=>'0', g4a=>'0');
  lcc_1c21 : ic_74s283 port map(s1    => lca1, b1 => gnd, a1 => lc1, s0 => lca0, a0 => lc0, b0 => internal25, c0 => lcinc, c4 => lcry3, s3 => lca3, b3 => gnd, a3 => lc3, s2 => lca2, a2 => lc2, b2 => gnd);
  lcc_1c27 : ic_25s09 port map(sel    => \-destlc\, aq => lc3, a0 => ob3, a1 => lca3, b1 => lca2, b0 => ob2, bq => lc2, clk => clk2a, cq => lc1, c0 => ob1, c1 => lca1, d1 => lca0, d0 => ob0, dq => lc0);
  lcc_1e07 : ic_74s08 port map(g4q    => lc0b, g4a => \lc_byte_mode\, g4b => lc0, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3a => '0', g3b => '0');
  lcc_2e05 : ic_74s86 port map(g1a    => \inst_in_left_half\, g1b => \-ir4\, g1y=>\-sh4\, g2a=>lc1, g2b=>lc0b, g2y=>internal27, g3y=>\-sh3\, g3a=>\-ir3\, g3b=>\inst_in_2nd_or_4th_quarter\, g4a=>'0', g4b=>'0');
  lcc_2e30 : ic_74s02 port map(g3b    => \-lc_modifies_mrot\, g3a => internal27, g3q_n => \inst_in_left_half\, g4b=>\-lc_modifies_mrot\, g4a=>lc0, g4q_n=>internal26, g1a=>'0', g1b=>'0', g2a=>'0', g2b=>'0');
  lcc_3e05 : ic_74s08 port map(g1b    => internal26, g1a => \lc_byte_mode\, g1q => \inst_in_2nd_or_4th_quarter\, g2b=>'0', g2a=>'0', g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');
  lcc_3e07 : ic_74s00 port map(g3q_n  => internal28, g3b => spc14, g3a => \-srcspcpopreal\, g4q_n => \-ifetch\, g4a=>needfetch, g4b=>lcinc, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0');
  lcc_3e09 : ic_74s32 port map(g4y    => needfetch, g4a => \have_wrong_word\, g4b => \last_byte_in_word\, g1a=>'0', g1b=>'0', g2a=>'0', g2b=>'0', g3a=>'0', g3b=>'0');
  lcc_3e11 : ic_74s00 port map(g1b    => ir10, g1a => ir11, g1q_n => \-lc_modifies_mrot\, g2b => \-newlc\, g2a=>\-destlc\, g2q_n=>\have_wrong_word\, g3q_n=>\-newlc.in\, g3b=>\-lcinc\, g3a=>\have_wrong_word\, g4a=>'0', g4b=>'0');
  lcc_3e12 : ic_74s175 port map(clr_n => \-reset\, q0 => \-newlc\, q0_n=>newlc, d0=>\-newlc.in\, d1=>int, q1_n=>nc359, q1=>sintr, clk=>clk3c, q2=>\next.instrd\, q2_n=>nc360, d2=>\next.instr\, d3=>nc361, q3_n=>nc362, q3=>nc363);
  lcc_3e17 : ic_74s02 port map(g1q_n  => \next.instr\, g1a => \-spop\, g1b=>internal28, g2q_n=>\last_byte_in_word\, g2a=>lc1, g2b=>lc0b, g3b=>internal29, g3a=>\next.instrd\, g3q_n=>\-lcinc\, g4b=>'0', g4a=>'0');
  lcc_3e22 : ic_74s04 port map(g3a    => needfetch, g3q_n => \-needfetch\, g1a => '0', g2a => '0', g4a => '0', g5a => '0', g6a => '0');
  lcc_4d09 : ic_74s08 port map(g2b    => spc14, g2a => \-needfetch\, g2q => spcmung, g4q => internal29, g4a => ir24, g4b => irdisp, g1b => '0', g1a => '0', g3a => '0', g3b => '0');
  lcc_4e03 : ic_74s32 port map(g1a    => spcmung, g1b => spc1, g1y => spc1a, g4y => lcinc, g4a => \next.instrd\, g4b => internal29, g2a => '0', g2b => '0', g3a => '0', g3b => '0');

  --- The VMA and VMA Selector

  vma_1a06 : ic_74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma31\, bout3=>mf24, ain1=>\-vma30\, bout2=>mf25, ain2=>\-vma29\, bout1=>mf26, ain3=>\-vma28\, bout0=>mf27, bin0=>\-vma27\, aout3=>mf28, bin1=>\-vma26\, aout2=>mf29, bin2=>\-vma25\, aout1=>mf30, bin3=>\-vma24\, aout0=>mf31, benb_n=>\-vmadrive\);
  vma_1a10 : ic_74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma7\, bout3=>mf0, ain1=>\-vma6\, bout2=>mf1, ain2=>\-vma5\, bout1=>mf2, ain3=>\-vma4\, bout0=>mf3, bin0=>\-vma3\, aout3=>mf4, bin1=>\-vma2\, aout2=>mf5, bin2=>\-vma1\, aout1=>mf6, bin3=>\-vma0\, aout0=>mf7, benb_n=>\-vmadrive\);
  vma_1a12 : ic_74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma23\, bout3=>mf16, ain1=>\-vma22\, bout2=>mf17, ain2=>\-vma21\, bout1=>mf18, ain3=>\-vma20\, bout0=>mf19, bin0=>\-vma19\, aout3=>mf20, bin1=>\-vma18\, aout2=>mf21, bin2=>\-vma17\, aout1=>mf22, bin3=>\-vma16\, aout0=>mf23, benb_n=>\-vmadrive\);
  vma_1a14 : ic_74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma15\, bout3=>mf8, ain1=>\-vma14\, bout2=>mf9, ain2=>\-vma13\, bout1=>mf10, ain3=>\-vma12\, bout0=>mf11, bin0=>\-vma11\, aout3=>mf12, bin1=>\-vma10\, aout2=>mf13, bin2=>\-vma9\, aout1=>mf14, bin3=>\-vma8\, aout0=>mf15, benb_n=>\-vmadrive\);
  vma_1a18 : ic_74s00 port map(g4q_n   => \-vmadrive\, g4a => tse2, g4b => srcvma, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3b => '0', g3a => '0');
  vma_1b22 : ic_25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma24\, i0=>\-vmas24\, i1=>\-vmas25\, d1=>\-vma25\, i2=>\-vmas26\, d2=>\-vma26\, clk=>clk1a, d3=>\-vma27\, i3=>\-vmas27\, d4=>\-vma28\, i4=>\-vmas28\, i5=>\-vmas29\, d5=>\-vma29\);
  vma_1b23 : ic_25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma30\, i0=>\-vmas30\, i1=>\-vmas31\, d1=>\-vma31\, i2=>nc115, d2=>nc116, clk=>clk1a, d3=>nc117, i3=>nc118, d4=>nc119, i4=>nc120, i5=>nc121, d5=>nc122);
  vma_1c22 : ic_25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma0\, i0=>\-vmas0\, i1=>\-vmas1\, d1=>\-vma1\, i2=>\-vmas2\, d2=>\-vma2\, clk=>clk2a, d3=>\-vma3\, i3=>\-vmas3\, d4=>\-vma4\, i4=>\-vmas4\, i5=>\-vmas5\, d5=>\-vma5\);
  vma_1c24 : ic_25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma12\, i0=>\-vmas12\, i1=>\-vmas13\, d1=>\-vma13\, i2=>\-vmas14\, d2=>\-vma14\, clk=>clk2a, d3=>\-vma15\, i3=>\-vmas15\, d4=>\-vma16\, i4=>\-vmas16\, i5=>\-vmas17\, d5=>\-vma17\);
  vma_1c25 : ic_25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma18\, i0=>\-vmas18\, i1=>\-vmas19\, d1=>\-vma19\, i2=>\-vmas20\, d2=>\-vma20\, clk=>clk2a, d3=>\-vma21\, i3=>\-vmas21\, d4=>\-vma22\, i4=>\-vmas22\, i5=>\-vmas23\, d5=>\-vma23\);
  vma_1d25 : ic_25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma6\, i0=>\-vmas6\, i1=>\-vmas7\, d1=>\-vma7\, i2=>\-vmas8\, d2=>\-vma8\, clk=>clk2c, d3=>\-vma9\, i3=>\-vmas9\, d4=>\-vma10\, i4=>\-vmas10\, i5=>\-vmas11\, d5=>\-vma11\);
  vma_2a05 : ic_74s04 port map(g3a     => \-srcvma\, g3q_n => srcvma, g1a => '0', g2a => '0', g4a => '0', g5a => '0', g6a => '0');

  vmas_1a27 : ic_74s258 port map(sel => vmasela, d0 => lc22, d1 => ob20, dy => \-vmas20\, c0 => lc23, c1 => ob21, cy => \-vmas21\, by=>\-vmas22\, b1=>ob22, b0=>lc24, ay=>\-vmas23\, a1=>ob23, a0=>lc25, enb_n=>gnd);
  vmas_1a29 : ic_74s258 port map(sel => vmasela, d0 => gnd, d1 => ob28, dy => \-vmas28\, c0 => gnd, c1 => ob29, cy => \-vmas29\, by=>\-vmas30\, b1=>ob30, b0=>gnd, ay=>\-vmas31\, a1=>ob31, a0=>gnd, enb_n=>gnd);
  vmas_1b26 : ic_74s258 port map(sel => vmaselb, d0 => lc14, d1 => ob12, dy => \-vmas12\, c0 => lc15, c1 => ob13, cy => \-vmas13\, by=>\-vmas14\, b1=>ob14, b0=>lc16, ay=>\-vmas15\, a1=>ob15, a0=>lc17, enb_n=>gnd);
  vmas_1b29 : ic_74s258 port map(sel => vmasela, d0 => lc18, d1 => ob16, dy => \-vmas16\, c0 => lc19, c1 => ob17, cy => \-vmas17\, by=>\-vmas18\, b1=>ob18, b0=>lc20, ay=>\-vmas19\, a1=>ob19, a0=>lc21, enb_n=>gnd);
  vmas_1c16 : ic_74s258 port map(sel => \-memstart\, d0 => \-vma12\, d1=>\-md12\, dy=>mapi12, c0=>\-vma13\, c1=>\-md13\, cy=>mapi13, by=>mapi14, b1=>\-md14\, b0=>\-vma14\, ay=>mapi15, a1=>\-md15\, a0=>\-vma15\, enb_n=>gnd);
  vmas_1c18 : ic_74s258 port map(sel => \-memstart\, d0 => \-vma16\, d1=>\-md16\, dy=>mapi16, c0=>\-vma17\, c1=>\-md17\, cy=>mapi17, by=>mapi18, b1=>\-md18\, b0=>\-vma18\, ay=>mapi19, a1=>\-md19\, a0=>\-vma19\, enb_n=>gnd);
  vmas_1c20 : ic_74s258 port map(sel => \-memstart\, d0 => \-vma20\, d1=>\-md20\, dy=>mapi20, c0=>\-vma21\, c1=>\-md21\, cy=>mapi21, by=>mapi22, b1=>\-md22\, b0=>\-vma22\, ay=>mapi23, a1=>\-md23\, a0=>\-vma23\, enb_n=>gnd);
  vmas_1c28 : ic_74s258 port map(sel => vmaselb, d0 => lc2, d1 => ob0, dy => \-vmas0\, c0 => lc3, c1 => ob1, cy => \-vmas1\, by=>\-vmas2\, b1=>ob2, b0=>lc4, ay=>\-vmas3\, a1=>ob3, a0=>lc5, enb_n=>gnd);
  vmas_1d19 : ic_74s258 port map(sel => \-memstart\, d0 => \-vma8\, d1=>\-md8\, dy=>mapi8, c0=>\-vma9\, c1=>\-md9\, cy=>mapi9, by=>mapi10, b1=>\-md10\, b0=>\-vma10\, ay=>mapi11, a1=>\-md11\, a0=>\-vma11\, enb_n=>gnd);
  vmas_1d30 : ic_74s258 port map(sel => vmaselb, d0 => lc10, d1 => ob8, dy => \-vmas8\, c0 => lc11, c1 => ob9, cy => \-vmas9\, by=>\-vmas10\, b1=>ob10, b0=>lc12, ay=>\-vmas11\, a1=>ob11, a0=>lc13, enb_n=>gnd);
  vmas_2b01 : ic_74s258 port map(sel => vmaselb, d0 => lc6, d1 => ob4, dy => \-vmas4\, c0 => lc7, c1 => ob5, cy => \-vmas5\, by=>\-vmas6\, b1=>ob6, b0=>lc8, ay=>\-vmas7\, a1=>ob7, a0=>lc9, enb_n=>gnd);
  vmas_2b04 : ic_74s258 port map(sel => vmasela, d0 => gnd, d1 => ob24, dy => \-vmas24\, c0 => gnd, c1 => ob25, cy => \-vmas25\, by=>\-vmas26\, b1=>ob26, b0=>gnd, ay=>\-vmas27\, a1=>ob27, a0=>gnd, enb_n=>gnd);

  --- The MD and the MD Selector

  md_1a02 : ic_74s240 port map(aenb_n => \-mddrive\, ain0 => \-md31\, bout3=>mf24, ain1=>\-md30\, bout2=>mf25, ain2=>\-md29\, bout1=>mf26, ain3=>\-md28\, bout0=>mf27, bin0=>\-md27\, aout3=>mf28, bin1=>\-md26\, aout2=>mf29, bin2=>\-md25\, aout1=>mf30, bin3=>\-md24\, aout0=>mf31, benb_n=>\-mddrive\);
  md_1a04 : ic_74s240 port map(aenb_n => \-mddrive\, ain0 => \-md23\, bout3=>mf16, ain1=>\-md22\, bout2=>mf17, ain2=>\-md21\, bout1=>mf18, ain3=>\-md20\, bout0=>mf19, bin0=>\-md19\, aout3=>mf20, bin1=>\-md18\, aout2=>mf21, bin2=>\-md17\, aout1=>mf22, bin3=>\-md16\, aout0=>mf23, benb_n=>\-mddrive\);
  md_1a05 : ic_74s240 port map(aenb_n => \-mddrive\, ain0 => \-md7\, bout3=>mf0, ain1=>\-md6\, bout2=>mf1, ain2=>\-md5\, bout1=>mf2, ain3=>\-md4\, bout0=>mf3, bin0=>\-md3\, aout3=>mf4, bin1=>\-md2\, aout2=>mf5, bin2=>\-md1\, aout1=>mf6, bin3=>\-md0\, aout0=>mf7, benb_n=>\-mddrive\);
  md_1a08 : ic_74s00 port map(g2b     => srcmd, g2a => tse2, g2q_n => \-mddrive\, g1b => '0', g1a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  md_1a09 : ic_74s240 port map(aenb_n => \-mddrive\, ain0 => \-md15\, bout3=>mf8, ain1=>\-md14\, bout2=>mf9, ain2=>\-md13\, bout1=>mf10, ain3=>\-md12\, bout0=>mf11, bin0=>\-md11\, aout3=>mf12, bin1=>\-md10\, aout2=>mf13, bin2=>\-md9\, aout1=>mf14, bin3=>\-md8\, aout0=>mf15, benb_n=>\-mddrive\);
  md_1b16 : ic_74s374 port map(oenb_n => gnd, o0 => \-md31\, i0 => \-mds31\, i1=>\-mds30\, o1=>\-md30\, o2=>\-md29\, i2=>\-mds29\, i3=>\-mds28\, o3=>\-md28\, clk=>mdclk, o4=>\-md27\, i4=>\-mds27\, i5=>\-mds26\, o5=>\-md26\, o6=>\-md25\, i6=>\-mds25\, i7=>\-mds24\, o7=>\-md24\);
  md_1c17 : ic_74s374 port map(oenb_n => gnd, o0 => \-md7\, i0 => \-mds7\, i1=>\-mds6\, o1=>\-md6\, o2=>\-md5\, i2=>\-mds5\, i3=>\-mds4\, o3=>\-md4\, clk=>mdclk, o4=>\-md3\, i4=>\-mds3\, i5=>\-mds2\, o5=>\-md2\, o6=>\-md1\, i6=>\-mds1\, i7=>\-mds0\, o7=>\-md0\);
  md_1c19 : ic_74s374 port map(oenb_n => gnd, o0 => \-md23\, i0 => \-mds23\, i1=>\-mds22\, o1=>\-md22\, o2=>\-md21\, i2=>\-mds21\, i3=>\-mds20\, o3=>\-md20\, clk=>mdclk, o4=>\-md19\, i4=>\-mds19\, i5=>\-mds18\, o5=>\-md18\, o6=>\-md17\, i6=>\-mds17\, i7=>\-mds16\, o7=>\-md16\);
  md_1d16 : ic_74s51 port map(g2a     => destmdr, g2b => \-clk2c\, g2c => loadmd, g2d => loadmd, g2y => mdclk, g1a => '0', g1c => '0', g1d => '0', g1b => '0');
  md_1d18 : ic_74s04 port map(g4q     => loadmd, g4a => \-loadmd\, g5q_n => destmdr, g5a => \-destmdr\, g1a=>'0', g2a=>'0', g3a=>'0', g6a=>'0');
  md_1d20 : ic_74s374 port map(oenb_n => gnd, o0 => \-md15\, i0 => \-mds15\, i1=>\-mds14\, o1=>\-md14\, o2=>\-md13\, i2=>\-mds13\, i3=>\-mds12\, o3=>\-md12\, clk=>mdclk, o4=>\-md11\, i4=>\-mds11\, i5=>\-mds10\, o5=>\-md10\, o6=>\-md9\, i6=>\-mds9\, i7=>\-mds8\, o7=>\-md8\);
  md_1e07 : ic_74s08 port map(g3q     => mdgetspar, g3a => \-destmdr\, g3b => \-ignpar\, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0', g4a=>'0', g4b=>'0');
  md_1e19 : ic_74s374 port map(oenb_n => gnd, o0 => nc322, i0 => nc323, i1 => nc324, o1 => nc325, o2 => nc326, i2 => nc327, i3 => nc328, o3 => nc329, clk => mdclk, o4 => nc330, i4 => nc331, i5 => nc332, o5 => nc333, o6 => mdhaspar, i6 => mdgetspar, i7 => \mempar_in\, o7 => mdpar);
  md_2a05 : ic_74s04 port map(g2a     => \-srcmd\, g2q_n => srcmd, g1a => '0', g3a => '0', g4a => '0', g5a => '0', g6a => '0');

  mds_1a11 : ic_74s240 port map(aenb_n => \-memdrive.a\, ain0 => \-md31\, bout3=>mem24, ain1=>\-md30\, bout2=>mem25, ain2=>\-md29\, bout1=>mem26, ain3=>\-md28\, bout0=>mem27, bin0=>\-md27\, aout3=>mem28, bin1=>\-md26\, aout2=>mem29, bin2=>\-md25\, aout1=>mem30, bin3=>\-md24\, aout0=>mem31, benb_n=>\-memdrive.b\);
  mds_1a15 : ic_74s240 port map(aenb_n => \-memdrive.a\, ain0 => \-md7\, bout3=>mem0, ain1=>\-md6\, bout2=>mem1, ain2=>\-md5\, bout1=>mem2, ain3=>\-md4\, bout0=>mem3, bin0=>\-md3\, aout3=>mem4, bin1=>\-md2\, aout2=>mem5, bin2=>\-md1\, aout1=>mem6, bin3=>\-md0\, aout0=>mem7, benb_n=>\-memdrive.b\);
  mds_1a17 : ic_74s240 port map(aenb_n => \-memdrive.a\, ain0 => \-md23\, bout3=>mem16, ain1=>\-md22\, bout2=>mem17, ain2=>\-md21\, bout1=>mem18, ain3=>\-md20\, bout0=>mem19, bin0=>\-md19\, aout3=>mem20, bin1=>\-md18\, aout2=>mem21, bin2=>\-md17\, aout1=>mem22, bin3=>\-md16\, aout0=>mem23, benb_n=>\-memdrive.b\);
  mds_1a19 : ic_74s240 port map(aenb_n => \-memdrive.a\, ain0 => \-md15\, bout3=>mem8, ain1=>\-md14\, bout2=>mem9, ain2=>\-md13\, bout1=>mem10, ain3=>\-md12\, bout0=>mem11, bin0=>\-md11\, aout3=>mem12, bin1=>\-md10\, aout2=>mem13, bin2=>\-md9\, aout1=>mem14, bin3=>\-md8\, aout0=>mem15, benb_n=>\-memdrive.b\);
  mds_1a28 : ic_74s258 port map(sel    => mdsela, d0 => mem20, d1 => ob20, dy => \-mds20\, c0 => mem21, c1 => ob21, cy => \-mds21\, by=>\-mds22\, b1=>ob22, b0=>mem22, ay=>\-mds23\, a1=>ob23, a0=>mem23, enb_n=>gnd);
  mds_1a30 : ic_74s258 port map(sel    => mdsela, d0 => mem28, d1 => ob28, dy => \-mds28\, c0 => mem29, c1 => ob29, cy => \-mds29\, by=>\-mds30\, b1=>ob30, b0=>mem30, ay=>\-mds31\, a1=>ob31, a0=>mem31, enb_n=>gnd);
  mds_1b05 : ic_74s240 port map(aenb_n => \-memdrive.a\, ain0 => nc308, bout3 => nc309, ain1 => nc310, bout2 => nc311, ain2 => nc312, bout1 => nc313, ain3 => mdparodd, bout0 => nc314, bin0 => nc315, aout3 => \mempar_out\, bin1=>nc316, aout2=>nc317, bin2=>nc318, aout1=>nc319, bin3=>nc320, aout0=>nc321, benb_n=>hi11);
  mds_1b27 : ic_74s258 port map(sel    => mdselb, d0 => mem12, d1 => ob12, dy => \-mds12\, c0 => mem13, c1 => ob13, cy => \-mds13\, by=>\-mds14\, b1=>ob14, b0=>mem14, ay=>\-mds15\, a1=>ob15, a0=>mem15, enb_n=>gnd);
  mds_1b30 : ic_74s258 port map(sel    => mdsela, d0 => mem16, d1 => ob16, dy => \-mds16\, c0 => mem17, c1 => ob17, cy => \-mds17\, by=>\-mds18\, b1=>ob18, b0=>mem18, ay=>\-mds19\, a1=>ob19, a0=>mem19, enb_n=>gnd);
  mds_1c26 : ic_74s258 port map(sel    => mdselb, d0 => mem8, d1 => ob8, dy => \-mds8\, c0 => mem9, c1 => ob9, cy => \-mds9\, by=>\-mds10\, b1=>ob10, b0=>mem10, ay=>\-mds11\, a1=>ob11, a0=>mem11, enb_n=>gnd);
  mds_1c29 : ic_74s258 port map(sel    => mdselb, d0 => mem0, d1 => ob0, dy => \-mds0\, c0 => mem1, c1 => ob1, cy => \-mds1\, by=>\-mds2\, b1=>ob2, b0=>mem2, ay=>\-mds3\, a1=>ob3, a0=>mem3, enb_n=>gnd);
  mds_2b02 : ic_74s258 port map(sel    => mdselb, d0 => mem4, d1 => ob4, dy => \-mds4\, c0 => mem5, c1 => ob5, cy => \-mds5\, by=>\-mds6\, b1=>ob6, b0=>mem6, ay=>\-mds7\, a1=>ob7, a0=>mem7, enb_n=>gnd);
  mds_2b05 : ic_74s258 port map(sel    => mdsela, d0 => mem24, d1 => ob24, dy => \-mds24\, c0 => mem25, c1 => ob25, cy => \-mds25\, by=>\-mds26\, b1=>ob26, b0=>mem26, ay=>\-mds27\, a1=>ob27, a0=>mem27, enb_n=>gnd);

  --- First and Second Level Maps

  vmem0_1c01 : ic_74s280 port map(i0   => \-vmap0\, i1 => \-vmap1\, i2=>\-vmap2\, even=>nc113, odd=>internal14, i3=>\-vmap3\, i4=>\-vmap4\, i5=>vpari, i6=>gnd, i7=>gnd, i8=>gnd);
  vmem0_1c02 : ic_74s280 port map(i0   => \-vma27\, i1 => \-vma28\, i2=>\-vma29\, even=>vm0pari, odd=>nc114, i3=>\-vma30\, i4=>\-vma31\, i5=>gnd, i6=>gnd, i7=>gnd, i8=>gnd);
  vmem0_1c06 : ic_93425a port map(ce_n => \-mapi23\, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap2\, a5=>mapi17, a6=>mapi16, a7=>mapi15, a8=>mapi14, a9=>mapi13, we_n=>\-vm0wpb\, di=>\-vma29\);
  vmem0_1c07 : ic_93425a port map(ce_n => mapi23, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap0\, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpa\, di=>\-vma27\);
  vmem0_1c08 : ic_93425a port map(ce_n => mapi23, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap1\, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpa\, di=>\-vma28\);
  vmem0_1c09 : ic_93425a port map(ce_n => mapi23, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap2\, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpa\, di=>\-vma29\);
  vmem0_1c11 : ic_93425a port map(ce_n => \-mapi23\, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap3\, a5=>mapi17, a6=>mapi16, a7=>mapi15, a8=>mapi14, a9=>mapi13, we_n=>\-vm0wpb\, di=>\-vma30\);
  vmem0_1c12 : ic_93425a port map(ce_n => \-mapi23\, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap4\, a5=>mapi17, a6=>mapi16, a7=>mapi15, a8=>mapi14, a9=>mapi13, we_n=>\-vm0wpb\, di=>\-vma31\);
  vmem0_1c13 : ic_93425a port map(ce_n => mapi23, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap3\, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpa\, di=>\-vma30\);
  vmem0_1c14 : ic_93425a port map(ce_n => mapi23, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap4\, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpa\, di=>\-vma31\);
  vmem0_1d04 : ic_93425a port map(ce_n => \-mapi23\, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => vpari, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpb\, di=>vm0pari);
  vmem0_1d05 : ic_93425a port map(ce_n => mapi23, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => vpari, a5 => mapi17, a6 => mapi16, a7 => mapi15, a8 => mapi14, a9 => mapi13, we_n => \-vm0wpa\, di => vm0pari);
  vmem0_1d09 : ic_93425a port map(ce_n => \-mapi23\, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap0\, a5=>mapi17, a6=>mapi16, a7=>mapi15, a8=>mapi14, a9=>mapi13, we_n=>\-vm0wpb\, di=>\-vma27\);
  vmem0_1d10 : ic_93425a port map(ce_n => \-mapi23\, a0 => mapi22, a1 => mapi21, a2 => mapi20, a3 => mapi19, a4 => mapi18, do => \-vmap1\, a5=>mapi17, a6=>mapi16, a7=>mapi15, a8=>mapi14, a9=>mapi13, we_n=>\-vm0wpb\, di=>\-vma28\);
  vmem0_1d18 : ic_74s04 port map(g1a   => mapi23, g1q_n => \-mapi23\, g2a => '0', g3a => '0', g4a => '0', g5a => '0', g6a => '0');
  vmem0_1d27 : ic_74s02 port map(g4b   => memstart, g4a => srcmap, g4q_n => \-use.map\, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g3b => '0', g3a => '0');
  vmem0_1e26 : ic_74s32 port map(g1a   => \-use.map\, g1b => internal14, g1y => v0parok, g2a => \-use.map\, g2b=>vmoparodd, g2y=>vmoparok, g3a=>'0', g3b=>'0', g4a=>'0', g4b=>'0');

  vmem1_1c03 : ic_93s48 port map(i6      => \-vma17\, i5 => \-vma18\, i4=>\-vma19\, i3=>\-vma20\, i2=>\-vma21\, i1=>\-vma22\, i0=>\-vma23\, po=>vm1mpar, pe=>nc109, i11=>\-vma12\, i10=>\-vma13\, i9=>\-vma14\, i8=>\-vma15\, i7=>\-vma16\);
  vmem1_1c04 : ic_93s48 port map(i6      => \-vma5\, i5 => \-vma6\, i4=>\-vma7\, i3=>\-vma8\, i2=>\-vma9\, i1=>\-vma10\, i0=>\-vma11\, po=>nc110, pe=>\-vm1lpar\, i11=>\-vma0\, i10=>\-vma1\, i9=>\-vma2\, i8=>\-vma3\, i7=>\-vma4\);
  vmem1_1d01 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo10\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma10\);
  vmem1_1d02 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo4\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma4\);
  vmem1_1d06 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo2\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma2\);
  vmem1_1d08 : ic_74s240 port map(aenb_n => gnd, ain0 => mapi10, bout3 => vmap0a, ain1 => mapi9, bout2 => vmap1a, ain2 => mapi8, bout1 => vmap2a, ain3 => \-vmap4\, bout0 => vmap3a, bin0 => \-vmap3\, aout3=>vmap4a, bin1=>\-vmap2\, aout2=>\-mapi8a\, bin2=>\-vmap1\, aout1=>\-mapi9a\, bin3=>\-vmap0\, aout0=>\-mapi10a\, benb_n=>gnd);
  vmem1_1d11 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo0\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma0\);
  vmem1_1d12 : ic_74s86 port map(g1a     => vm1mpar, g1b => \-vm1lpar\, g1y => vm1pari, g2a => '0', g2b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  vmem1_1d13 : ic_74s240 port map(aenb_n => gnd, ain0 => mapi12, bout3 => \-mapi11a\, ain1 => mapi11, bout2 => \-mapi12a\, ain2=>mapi10, bout1=>nc111, ain3=>mapi9, bout0=>\-mapi8b\, bin0=>mapi8, aout3=>\-mapi9b\, bin1=>nc112, aout2=>\-mapi10b\, bin2=>mapi12, aout1=>\-mapi11b\, bin3=>mapi11, aout0=>\-mapi12b\, benb_n=>gnd);
  vmem1_1e04 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo11\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma11\);
  vmem1_1e05 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo5\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma5\);
  vmem1_1e08 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo9\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma9\);
  vmem1_1e09 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo3\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma3\);
  vmem1_1e10 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo8\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma8\);
  vmem1_1e13 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo7\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma7\);
  vmem1_1e14 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo1\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma1\);
  vmem1_1e15 : ic_93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo6\, a5 => \-mapi12a\, a6=>\-mapi11a\, a7=>\-mapi10a\, a8=>\-mapi9a\, a9=>\-mapi8a\, we_n=>\-vm1wpa\, di=>\-vma6\);

  vmem2_1b01 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo20\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma20\);
  vmem2_1b02 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo21\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma21\);
  vmem2_1b03 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo22\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma22\);
  vmem2_1b04 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo23\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma23\);
  vmem2_1b06 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo16\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma16\);
  vmem2_1b07 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo17\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma17\);
  vmem2_1b08 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo18\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma18\);
  vmem2_1b09 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo19\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma19\);
  vmem2_1b11 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo12\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma12\);
  vmem2_1b12 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo13\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma13\);
  vmem2_1b13 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo14\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma14\);
  vmem2_1b14 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => \-vmo15\, a5 => \-mapi12b\, a6=>\-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>\-vma15\);
  vmem2_1b17 : ic_93s48 port map(i6      => \-vmo17\, i5 => \-vmo18\, i4=>\-vmo19\, i3=>\-vmo20\, i2=>\-vmo21\, i1=>\-vmo22\, i0=>\-vmo23\, po=>vmoparm, pe=>nc107, i11=>\-vmo12\, i10=>\-vmo13\, i9=>\-vmo14\, i8=>\-vmo15\, i7=>\-vmo16\);
  vmem2_1c05 : ic_93425a port map(ce_n   => gnd, a0 => vmap4b, a1 => vmap3b, a2 => vmap2b, a3 => vmap1b, a4 => vmap0b, do => vmopar, a5 => \-mapi12b\, a6 => \-mapi11b\, a7=>\-mapi10b\, a8=>\-mapi9b\, a9=>\-mapi8b\, we_n=>\-vm1wpb\, di=>vm1pari);
  vmem2_1c10 : ic_74s240 port map(aenb_n => gnd, ain0 => nc101, bout3 => vmap0b, ain1 => nc102, bout2 => vmap1b, ain2 => nc103, bout1 => vmap2b, ain3 => \-vmap4\, bout0 => vmap3b, bin0 => \-vmap3\, aout3=>vmap4b, bin1=>\-vmap2\, aout2=>nc104, bin2=>\-vmap1\, aout1=>nc105, bin3=>\-vmap0\, aout0=>nc106, benb_n=>gnd);
  vmem2_1d03 : ic_93s48 port map(i6      => \-vmo5\, i5 => \-vmo6\, i4=>\-vmo7\, i3=>\-vmo8\, i2=>\-vmo9\, i1=>\-vmo10\, i0=>\-vmo11\, po=>vmoparl, pe=>nc108, i11=>\-vmo0\, i10=>\-vmo1\, i9=>\-vmo2\, i8=>\-vmo3\, i7=>\-vmo4\);
  vmem2_1d12 : ic_74s86 port map(g2a     => vmoparm, g2b => vmoparl, g2y => vmoparck, g3y => vmoparodd, g3a => vmopar, g3b => vmoparck, g1a => '0', g1b => '0', g4a => '0', g4b => '0');

  vmemdr_1a01 : ic_74s240 port map(aenb_n => \-mapdrive\, ain0 => \-pfw\, bout3=>mf24, ain1=>\-pfr\, bout2=>mf25, ain2=>hi12, bout1=>mf26, ain3=>\-vmap4\, bout0=>mf27, bin0=>\-vmap3\, aout3=>mf28, bin1=>\-vmap2\, aout2=>mf29, bin2=>\-vmap1\, aout1=>mf30, bin3=>\-vmap0\, aout0=>mf31, benb_n=>\-mapdrive\);
  vmemdr_1a03 : ic_74s240 port map(aenb_n => \-mapdrive\, ain0 => \-vmo15\, bout3=>mf8, ain1=>\-vmo14\, bout2=>mf9, ain2=>\-vmo13\, bout1=>mf10, ain3=>\-vmo12\, bout0=>mf11, bin0=>\-vmo11\, aout3=>mf12, bin1=>\-vmo10\, aout2=>mf13, bin2=>\-vmo9\, aout1=>mf14, bin3=>\-vmo8\, aout0=>mf15, benb_n=>\-mapdrive\);
  vmemdr_1a07 : ic_74s240 port map(aenb_n => \-mapdrive\, ain0 => \-vmo23\, bout3=>mf16, ain1=>\-vmo22\, bout2=>mf17, ain2=>\-vmo21\, bout1=>mf18, ain3=>\-vmo20\, bout0=>mf19, bin0=>\-vmo19\, aout3=>mf20, bin1=>\-vmo18\, aout2=>mf21, bin2=>\-vmo17\, aout1=>mf22, bin3=>\-vmo16\, aout0=>mf23, benb_n=>\-mapdrive\);
  vmemdr_1a08 : ic_74s00 port map(g1b     => tse1a, g1a => srcmap, g1q_n => \-mapdrive\, g2b => '0', g2a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  vmemdr_1a13 : ic_74s240 port map(aenb_n => \-mapdrive\, ain0 => \-vmo7\, bout3=>mf0, ain1=>\-vmo6\, bout2=>mf1, ain2=>\-vmo5\, bout1=>mf2, ain3=>\-vmo4\, bout0=>mf3, bin0=>\-vmo3\, aout3=>mf4, bin1=>\-vmo2\, aout2=>mf5, bin2=>\-vmo1\, aout1=>mf6, bin3=>\-vmo0\, aout0=>mf7, benb_n=>\-mapdrive\);
  vmemdr_1d14 : ic_74s373 port map(oenb_n => gnd, o0 => \-lvmo23\, i0 => \-vmo23\, i1=>\-vmo22\, o1=>\-lvmo22\, o2=>\-pma21\, i2=>\-vmo13\, i3=>\-vmo12\, o3=>\-pma20\, hold_n=>memstart, o4=>\-pma19\, i4=>\-vmo11\, i5=>\-vmo10\, o5=>\-pma18\, o6=>\-pma17\, i6=>\-vmo9\, i7=>\-vmo8\, o7=>\-pma16\);
  vmemdr_1d15 : ic_74s373 port map(oenb_n => gnd, o0 => \-pma15\, i0 => \-vmo7\, i1=>\-vmo6\, o1=>\-pma14\, o2=>\-pma13\, i2=>\-vmo5\, i3=>\-vmo4\, o3=>\-pma12\, hold_n=>memstart, o4=>\-pma11\, i4=>\-vmo3\, i5=>\-vmo2\, o5=>\-pma10\, o6=>\-pma9\, i6=>\-vmo1\, i7=>\-vmo0\, o7=>\-pma8\);
  vmemdr_1e17 : ic_93s48 port map(i6      => \-vma6\, i5 => \-vma5\, i4=>\-vma4\, i3=>\-vma3\, i2=>\-vma2\, i1=>\-vma1\, i0=>\-vma0\, po=>internal13, pe=>nc100, i11=>\-pma11\, i10=>\-pma10\, i9=>\-pma9\, i8=>\-pma8\, i7=>\-vma7\);
  vmemdr_1e18 : ic_93s48 port map(i6      => \-pma18\, i5 => \-pma17\, i4=>\-pma16\, i3=>\-pma15\, i2=>\-pma14\, i1=>\-pma13\, i0=>\-pma12\, po=>\-adrpar\, pe=>nc99, i11=>internal13, i10=>gnd, i9=>\-pma21\, i8=>\-pma20\, i7=>\-pma19\);
  vmemdr_2a05 : ic_74s04 port map(g4q     => srcmap, g4a => \-srcmap\, g1a => '0', g2a => '0', g3a => '0', g5a => '0', g6a => '0');

  --- Memory Control Logic

  vctl1_1c23 : ic_74s175 port map(clr_n => \-reset\, q0 => nc126, q0_n => nc127, d0 => nc128, d1 => internal15, q1_n => rdcyc, q1 => wrcyc, clk => clk2a, q2 => nc129, q2_n => nc130, d2 => nc131, d3 => wmap, q3_n => \-wmapd\, q3=>wmapd);
  vctl1_1d16 : ic_74s51 port map(g1a    => rdcyc, g1y => internal15, g1c => memprepare, g1d => \-memwr\, g1b => \-memprepare\, g2a=>'0', g2b=>'0', g2c=>'0', g2d=>'0');
  vctl1_1d17 : ic_74s00 port map(g1b    => \-lvmo22\, g1a => wrcyc, g1q_n => \-pfw\, g2b=>\-pfr\, g2a=>\-pfw\, g2q_n=>\-vmaok\, g3b=>'0', g3a=>'0', g4a=>'0', g4b=>'0');
  vctl1_1d21 : ic_74s74 port map(g1r_n  => \-mfinishd\, g1d => memrq, g1clk => mclk1a, g1s_n => hi11, g1q => mbusy, g1q_n => nc139, g2q_n => nc140, g2q => \rd.in.progress\, g2s_n=>hi11, g2clk=>mclk1a, g2d=>\set.rd.in.progress\, g2r_n=>\-rdfinish\);
  vctl1_1d22 : ic_td250 port map(input  => internal16, o_100ns => \-rdfinish\, o_200ns => nc132, o_250ns => nc133, o_150ns => nc134, o_50ns => nc135);
  vctl1_1d23 : ic_td50 port map(input   => \-mfinish\, o_20ns => nc136, o_40ns => internal16, o_50ns => nc137, o_30ns => \-mfinishd\, o_10ns=>nc138);
  vctl1_1d27 : ic_74s02 port map(g3b    => clk2c, g3a => \-memop\, g3q_n => memprepare, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4b => '0', g4a => '0');
  vctl1_1d28 : ic_74s08 port map(g4q    => \-mfinish\, g4a => \-reset\, g4b=>\-memack\, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0', g3a=>'0', g3b=>'0');
  vctl1_1e16 : ic_74s11 port map(g2a    => \-memrd\, g2b => \-memwr\, g2c=>\-ifetch\, g2y_n=>\-memop\, g1a=>'0', g1b=>'0', g3a=>'0', g3b=>'0', g3c=>'0', g1c=>'0');
  vctl1_1e20 : ic_74s175 port map(clr_n => \-reset\, q0 => memstart, q0_n => \-memstart\, d0=>memprepare, d1=>memrq, q1_n=>\-mbusy.sync\, q1=>\mbusy.sync\, clk=>mclk1a, q2=>nc141, q2_n=>nc142, d2=>nc143, d3=>nc144, q3_n=>nc145, q3=>nc146);
  vctl1_1e25 : ic_9s42_1 port map(g1a1  => mbusy, g1b1 => hi11, g2a1 => memstart, g2b1 => \-pfr\, g2c1 => \-pfw\, g2d1=>hi11, out1=>memrq, out2=>\set.rd.in.progress\, g2d2=>hi11, g2c2=>rdcyc, g2b2=>\-pfr\, g2a2=>memstart, g1b2=>hi11, g1a2=>\rd.in.progress\);
  vctl1_3f16 : ic_74s64 port map(d4     => hi4, b2 => \mbusy.sync\, a2 => destmem, c3 => \-memgrant\, b3=>mbusy, a3=>\use.md\, \out\=>\-wait\, a1=>gnd, b1=>gnd, c4=>\mbusy.sync\, b4=>needfetch, a4=>lcinc);
  vctl1_3f17 : ic_74s10 port map(g1a    => \rd.in.progress\, g1b => \use.md\, g1y_n=>\-hang\, g1c=>\-clk3g\, g2a=>'0', g2b=>'0', g2c=>'0', g3a=>'0', g3b=>'0', g3c=>'0');

  vctl2_1c15 : ic_74s02 port map(g1q_n => mapwr0d, g1a => \-wmapd\, g1b => \-vma26\, g2q_n=>mapwr1d, g2a=>\-wmapd\, g2b=>\-vma25\, g3b=>'0', g3a=>'0', g4b=>'0', g4a=>'0');
  vctl2_1d07 : ic_74s37 port map(g1a   => mapwr0d, g1b => wp1a, g1y => \-vm0wpa\, g2a => mapwr0d, g2b => wp1a, g2y => \-vm0wpb\, g3y=>\-vm1wpa\, g3a=>wp1b, g3b=>mapwr1d, g4y=>\-vm1wpb\, g4a=>wp1b, g4b=>mapwr1d);
  vctl2_1d26 : ic_74s04 port map(g1a   => nc123, g1q_n => nc124, g2a => \-lvmo23\, g2q_n => \-pfr\, g3a=>\-wmap\, g3q_n=>wmap, g4q=>\-memrq\, g4a=>memrq, g5q_n=>\-memprepare\, g5a=>memprepare, g6q_n=>destmem, g6a=>\-destmem\);
  vctl2_1d27 : ic_74s02 port map(g1q_n => mdsela, g1a => \-destmdr\, g1b => clk2c, g2q_n => mdselb, g2a => \-destmdr\, g2b=>clk2c, g3b=>'0', g3a=>'0', g4b=>'0', g4a=>'0');
  vctl2_1d28 : ic_74s08 port map(g1b   => \-destvma\, g1a => \-ifetch\, g1q=>\-vmaenb\, g2b=>\-ifetch\, g2a=>hi11, g2q=>vmasela, g3q=>vmaselb, g3a=>hi11, g3b=>\-ifetch\, g4a=>'0', g4b=>'0');
  vctl2_1e06 : ic_74s00 port map(g1b   => wrcyc, g1a => \lm_drive_enb\, g1q_n => \-memdrive.a\, g2b=>wrcyc, g2a=>\lm_drive_enb\, g2q_n=>\-memdrive.b\, g3b=>'0', g3a=>'0', g4a=>'0', g4b=>'0');
  vctl2_3d04 : ic_74s139 port map(g2y3 => \-wmap\, g2y2 => \-memwr\, g2y1=>\-memrd\, g2y0=>nc125, b2=>ir20, a2=>ir19, g2=>\-destmem\, g1=>'0', a1=>'0', b1=>'0');
  vctl2_3f18 : ic_74s02 port map(g1q_n => \use.md\, g1a => \-srcmd\, g1b=>nopa, g2a=>'0', g2b=>'0', g3b=>'0', g3a=>'0', g4b=>'0', g4a=>'0');
  vctl2_3f19 : ic_74s04 port map(g5q_n => nopa, g5a => \-nopa\, g1a => '0', g2a => '0', g3a => '0', g4a => '0', g6a => '0');

  olord1_1a01 : ic_74s174 port map(clr_n => \-clock_reset_a\, q1 => nc84, d1 => nc85, d2 => nc86, q2 => nc87, d3 => speed1a, q3 => sspeed1, clk => speedclk, q4 => sspeed0, d4 => speed0a, q5 => speed1a, d5 => speed1, d6 => speed0, q6 => speed0a);
  olord1_1a04 : ic_74s174 port map(clr_n => \-reset\, q1 => speed0, d1 => spy0, d2 => spy1, q2 => speed1, d3 => spy2, q3 => errstop, clk => \-ldmode\, q4=>stathenb, d4=>spy3, q5=>trapenb, d5=>spy4, d6=>spy5, q6=>promdisable);
  olord1_1a08 : ic_74s175 port map(clr_n => \-reset\, q0 => nc92, q0_n => nc93, d0 => spy3, d1 => spy2, q1_n => \-opcinh\, q1=>opcinh, clk=>\-ldopc\, q2=>opcclk, q2_n=>\-opcclk\, d2=>spy1, d3=>spy0, q3_n=>\-lpc.hold\, q3=>\lpc.hold\);
  olord1_1a09 : ic_74s175 port map(clr_n => \-reset\, q0 => ldstat, q0_n => \-ldstat\, d0=>spy4, d1=>spy3, q1_n=>\-idebug\, q1=>idebug, clk=>\-ldclk\, q2=>nop11, q2_n=>\-nop11\, d2=>spy2, d3=>spy1, q3_n=>\-step\, q3=>step);
  olord1_1a10 : ic_74s174 port map(clr_n => \-clock_reset_a\, q1 => promdisabled, d1 => promdisable, d2 => sstep, q2 => ssdone, d3 => step, q3 => sstep, clk => mclk5a, q4 => srun, d4 => run, q5 => nc88, d5 => nc89, d6 => nc90, q6 => nc91);
  olord1_1a14 : ic_74s74 port map(g1r_n  => \-clock_reset_a\, g1d => spy0, g1clk => \-ldclk\, g1s_n=>\-boot\, g1q=>run, g1q_n=>\-run\, g2s_n=>'0', g2clk=>'0', g2d=>'0', g2r_n=>'0');
  olord1_1a15 : ic_9s42_1 port map(g1a1  => sstep, g1b1 => \-ssdone\, g2a1 => srun, g2b1 => \-errhalt\, g2c1=>\-wait\, g2d1=>\-stathalt\, out1=>machrun, g1a2=>'0', g1b2=>'0', g2a2=>'0', g2b2=>'0', g2c2=>'0', g2d2=>'0');
  olord1_1b10 : ic_74s04 port map(g2a    => ssdone, g2q_n => \-ssdone\, g5q_n => \stat.ovf\, g5a=>\-stc32\, g1a=>'0', g3a=>'0', g4a=>'0', g6a=>'0');
  olord1_1c01 : ic_7428 port map(g3a     => \-tpr60\, g3b => gnd, g3q_n => speedclk, g1a => '0', g1b => '0', g2a => '0', g4a => '0', g4b => '0', g2b => '0');
  olord1_1c09 : ic_74s00 port map(g3q_n  => \-stathalt\, g3b => stathenb, g3a => statstop, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  olord1_1c10 : ic_74s02 port map(g1q_n  => \-machruna\, g1a => gnd, g1b => machrun, g2a => '0', g2b => '0', g3b => '0', g3a => '0', g4b => '0', g4a => '0');
  olord1_1f10 : ic_74s04 port map(g4q    => \-machrun\, g4a => machrun, g1a => '0', g2a => '0', g3a => '0', g5a => '0', g6a => '0');

  olord2_1a02 : ic_74s133 port map(g       => \-ape\, f => \-mpe\, e=>\-pdlpe\, d=>\-dpe\, c=>\-ipe\, b=>\-spe\, a=>\-higherr\, q_n=>err, h=>\-mempe\, i=>\-v0pe\, j=>\-v1pe\, k=>\-halted\, l=>hi1, m=>hi1);
  olord2_1a03 : ic_74s374 port map(oenb_n  => gnd, o0 => \-ape\, i0 => aparok, i1 => mmemparok, o1 => \-mpe\, o2=>\-pdlpe\, i2=>pdlparok, i3=>dparok, o3=>\-dpe\, clk=>clk5a, o4=>\-ipe\, i4=>iparok, i5=>spcparok, o5=>\-spe\, o6=>\-higherr\, i6=>highok, i7=>memparok, o7=>\-mempe\);
  olord2_1a05 : ic_74s374 port map(oenb_n  => gnd, o0 => \-v0pe\, i0 => v0parok, i1 => vmoparok, o1 => \-v1pe\, o2=>statstop, i2=>\stat.ovf\, i3=>\-halt\, o3=>\-halted\, clk=>clk5a, o4=>nc76, i4=>nc77, i5=>nc78, o5=>nc79, o6=>nc80, i6=>nc81, i7=>nc82, o7=>nc83);
  olord2_1a06 : ic_74s37 port map(g1a      => \-mclk5\, g1b => \-mclk5\, g1y=>mclk5a, g2a=>\-clk5\, g2b=>\-clk5\, g2y=>clk5a, g3y=>\-reset\, g3a=>hi1, g3b=>reset, g4y=>\bus.power.reset_l\, g4a=>\power_reset_a\, g4b=>\power_reset_a\);
  olord2_1a07 : ic_74s02 port map(g1q_n    => highok, g1a => \-upperhighok\, g1b => \-lowerhighok\, g2q_n=>\-boot\, g2a=>internal5, g2b=>internal2, g3b=>\power_reset_a\, g3a=>\prog.bus.reset\, g3q_n=>\-bus.reset\, g4b=>'0', g4a=>'0');
  olord2_1a11 : ic_74s02 port map(g1q_n    => \-clock_reset_b\, g1a => \power_reset_a\, g1b=>internal1, g2q_n=>\-clock_reset_a\, g2a=>\power_reset_a\, g2b=>internal1, g3b=>gnd, g3a=>\-power_reset\, g3q_n=>\power_reset_a\, g4b=>'0', g4a=>'0');
  olord2_1a18 : ic_74ls109 port map(clr1_n => \-boot\, j1 => srun, k1_n => hi1, clk1 => mclk5a, pre1_n => \-clock_reset_a\, q1=>nc75, q1_n=>\boot.trap\, clr2_n=>'0', j2=>'0', k2_n=>'0', clk2=>'0', pre2_n=>'0');
  olord2_1a19 : ic_16dummy port map(dummy  => vcc);
  olord2_1a20 : ic_74ls14 port map(g1q_n   => internal4, g2a => \-boot1\, g2q_n => internal5, g3a => \-boot2\, g3q_n=>internal3, g4q=>\-power_reset\, g4a=>internal4, g1a=>'0', g5a=>'0', g6a=>'0');
  olord2_1b10 : ic_74s04 port map(g1a      => \-ldmode\, g1q_n => ldmode, g3a => mclk5, g3q_n => \-mclk5\, g4q=>\-clk5\, g4a=>clk5, g6q_n=>internal1, g6a=>\-busint.lm.reset\, g2a=>'0', g5a=>'0');
  olord2_1c07 : ic_74s00 port map(g4q_n    => \-lowerhighok\, g4a => hi2, g4b => hi1, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3b => '0', g3a => '0');
  olord2_1c08 : ic_74s10 port map(g3y_n    => reset, g3a => \-boot\, g3b => \-clock_reset_b\, g3c=>\-prog.reset\, g1a=>'0', g1b=>'0', g2a=>'0', g2b=>'0', g2c=>'0', g1c=>'0');
  olord2_1c09 : ic_74s00 port map(g2b      => ldmode, g2a => spy6, g2q_n => \-prog.reset\, g4q_n => \-errhalt\, g4a=>errstop, g4b=>err, g1b=>'0', g1a=>'0', g3b=>'0', g3a=>'0');
  olord2_1c18 : ic_74s32 port map(g3y      => internal2, g3a => internal3, g3b => \prog.boot\, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4a => '0', g4b => '0');
  olord2_1d10 : ic_74s08 port map(g2b      => ldmode, g2a => spy7, g2q => \prog.boot\, g1b => '0', g1a => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');

  --- Other

  stat_1b01 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr12, i1 => iwr13, i2 => iwr14, i3 => iwr15, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc12\, o3=>st15, o2=>st14, o1=>st13, o0=>st12, co_n=>\-stc16\);
  stat_1b02 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr16, i1 => iwr17, i2 => iwr18, i3 => iwr19, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc16\, o3=>st19, o2=>st18, o1=>st17, o0=>st16, co_n=>\-stc20\);
  stat_1b03 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr20, i1 => iwr21, i2 => iwr22, i3 => iwr23, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc20\, o3=>st23, o2=>st22, o1=>st21, o0=>st20, co_n=>\-stc24\);
  stat_1b04 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr24, i1 => iwr25, i2 => iwr26, i3 => iwr27, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc24\, o3=>st27, o2=>st26, o1=>st25, o0=>st24, co_n=>\-stc28\);
  stat_1b05 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr28, i1 => iwr29, i2 => iwr30, i3 => iwr31, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc28\, o3=>st31, o2=>st30, o1=>st29, o0=>st28, co_n=>\-stc32\);
  stat_1b06 : ic_74ls244 port map(aenb_n => \-spy.sth\, ain0 => st31, bout3 => spy8, ain1 => st30, bout2 => spy9, ain2 => st29, bout1 => spy10, ain3 => st28, bout0 => spy11, bin0 => st27, aout3 => spy12, bin1 => st26, aout2 => spy13, bin2 => st25, aout1 => spy14, bin3 => st24, aout0 => spy15, benb_n => \-spy.sth\);
  stat_1b07 : ic_74ls244 port map(aenb_n => \-spy.sth\, ain0 => st23, bout3 => spy0, ain1 => st22, bout2 => spy1, ain2 => st21, bout1 => spy2, ain3 => st20, bout0 => spy3, bin0 => st19, aout3 => spy4, bin1 => st18, aout2 => spy5, bin2 => st17, aout1 => spy6, bin3 => st16, aout0 => spy7, benb_n => \-spy.sth\);
  stat_1b08 : ic_74ls244 port map(aenb_n => \-spy.stl\, ain0 => st15, bout3 => spy8, ain1 => st14, bout2 => spy9, ain2 => st13, bout1 => spy10, ain3 => st12, bout0 => spy11, bin0 => st11, aout3 => spy12, bin1 => st10, aout2 => spy13, bin2 => st9, aout1 => spy14, bin3 => st8, aout0 => spy15, benb_n => \-spy.stl\);
  stat_1b09 : ic_74ls244 port map(aenb_n => \-spy.stl\, ain0 => st7, bout3 => spy0, ain1 => st6, bout2 => spy1, ain2 => st5, bout1 => spy2, ain3 => st4, bout0 => spy3, bin0 => st3, aout3 => spy4, bin1 => st2, aout2 => spy5, bin2 => st1, aout1 => spy6, bin3 => st0, aout0 => spy7, benb_n => \-spy.stl\);
  stat_1c03 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr0, i1 => iwr1, i2 => iwr2, i3 => iwr3, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-statbit\, o3=>st3, o2=>st2, o1=>st1, o0=>st0, co_n=>\-stc4\);
  stat_1c04 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr4, i1 => iwr5, i2 => iwr6, i3 => iwr7, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc4\, o3=>st7, o2=>st6, o1=>st5, o0=>st4, co_n=>\-stc8\);
  stat_1c05 : ic_74s169 port map(up_dn   => hi1, clk => clk5a, i0 => iwr8, i1 => iwr9, i2 => iwr10, i3 => iwr11, enb_p_n => gnd, load_n => \-ldstat\, enb_t_n => \-stc8\, o3=>st11, o2=>st10, o1=>st9, o0=>st8, co_n=>\-stc12\);

  opcs_1f06 : ic_9328 port map(clr_n  => hi2, aq_n => nc71, aq => opc13, asel => gnd, ai1 => nc72, ai0 => pc13, aclk => opcinha, comclk => opcclka, bclk => opcinha, bi0 => pc12, bi1 => nc73, bsel => gnd, bq => opc12, bq_n => nc74);
  opcs_1f07 : ic_9328 port map(clr_n  => hi2, aq_n => nc67, aq => opc11, asel => gnd, ai1 => nc68, ai0 => pc11, aclk => opcinha, comclk => opcclka, bclk => opcinha, bi0 => pc10, bi1 => nc69, bsel => gnd, bq => opc10, bq_n => nc70);
  opcs_1f08 : ic_9328 port map(clr_n  => hi2, aq_n => nc63, aq => opc9, asel => gnd, ai1 => nc64, ai0 => pc9, aclk => opcinha, comclk => opcclkc, bclk => opcinha, bi0 => pc8, bi1 => nc65, bsel => gnd, bq => opc8, bq_n => nc66);
  opcs_1f09 : ic_9328 port map(clr_n  => hi2, aq_n => nc59, aq => opc7, asel => gnd, ai1 => nc60, ai0 => pc7, aclk => opcinha, comclk => opcclkc, bclk => opcinha, bi0 => pc6, bi1 => nc61, bsel => gnd, bq => opc6, bq_n => nc62);
  opcs_1f10 : ic_74s04 port map(g1a   => \-opcinh\, g1q_n => opcinha, g2a => \-opcinh\, g2q_n=>opcinhb, g3a=>'0', g4a=>'0', g5a=>'0', g6a=>'0');
  opcs_1f11 : ic_9328 port map(clr_n  => hi2, aq_n => nc55, aq => opc5, asel => gnd, ai1 => nc56, ai0 => pc5, aclk => opcinhb, comclk => opcclkb, bclk => opcinhb, bi0 => pc4, bi1 => nc57, bsel => gnd, bq => opc4, bq_n => nc58);
  opcs_1f12 : ic_9328 port map(clr_n  => hi2, aq_n => nc51, aq => opc3, asel => gnd, ai1 => nc52, ai0 => pc3, aclk => opcinhb, comclk => opcclkb, bclk => opcinhb, bi0 => pc2, bi1 => nc53, bsel => gnd, bq => opc2, bq_n => nc54);
  opcs_1f13 : ic_9328 port map(clr_n  => hi2, aq_n => nc47, aq => opc1, asel => gnd, ai1 => nc48, ai0 => pc1, aclk => opcinhb, comclk => opcclkb, bclk => opcinhb, bi0 => pc0, bi1 => nc49, bsel => gnd, bq => opc0, bq_n => nc50);
  opcs_1f14 : ic_74s02 port map(g1q_n => opcclka, g1a => \-clk5\, g1b => opcclk, g2q_n => opcclkb, g2a => \-clk5\, g2b=>opcclk, g3b=>opcclk, g3a=>\-clk5\, g3q_n=>opcclkc, g4b=>'0', g4a=>'0');

  iwrpar_1b11 : ic_93s48 port map(i6 => iwr41, i5 => iwr42, i4 => iwr43, i3 => iwr44, i2 => iwr45, i1 => iwr46, i0 => iwr47, po => iwrp4, pe => nc98, i11 => iwr36, i10 => iwr37, i9 => iwr38, i8 => iwr39, i7 => iwr40);
  iwrpar_1b12 : ic_93s48 port map(i6 => iwr29, i5 => iwr30, i4 => iwr31, i3 => iwr32, i2 => iwr33, i1 => iwr34, i0 => iwr35, po => iwrp3, pe => nc97, i11 => iwr24, i10 => iwr25, i9 => iwr26, i8 => iwr27, i7 => iwr28);
  iwrpar_1b13 : ic_93s48 port map(i6 => iwr17, i5 => iwr18, i4 => iwr19, i3 => iwr20, i2 => iwr21, i1 => iwr22, i0 => iwr23, po => iwrp2, pe => nc96, i11 => iwr12, i10 => iwr13, i9 => iwr14, i8 => iwr15, i7 => iwr16);
  iwrpar_1b14 : ic_93s48 port map(i6 => iwr5, i5 => iwr6, i4 => iwr7, i3 => iwr8, i2 => iwr9, i1 => iwr10, i0 => iwr11, po => iwrp1, pe => nc95, i11 => iwr0, i10 => iwr1, i9 => iwr2, i8 => iwr3, i7 => iwr4);
  iwrpar_1b15 : ic_93s48 port map(i6 => gnd, i5 => gnd, i4 => gnd, i3 => gnd, i2 => gnd, i1 => gnd, i0 => gnd, po => nc94, pe => iwr48, i11 => iwrp1, i10 => iwrp2, i9 => iwrp3, i8 => iwrp4, i7 => gnd);

  trap_1d12 : ic_74s86 port map(g4y   => mdparerr, g4a => mdpareven, g4b => mdpar, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g3a => '0', g3b => '0');
  trap_1e28 : ic_93s48 port map(i6    => \-md5\, i5 => \-md6\, i4=>\-md7\, i3=>\-md8\, i2=>\-md9\, i1=>\-md10\, i0=>\-md11\, po=>mdparl, pe=>nc148, i11=>\-md0\, i10=>\-md1\, i9=>\-md2\, i8=>\-md3\, i7=>\-md4\);
  trap_1e29 : ic_93s48 port map(i6    => \-md17\, i5 => \-md18\, i4=>\-md19\, i3=>\-md20\, i2=>\-md21\, i1=>\-md22\, i0=>\-md23\, po=>mdparm, pe=>nc147, i11=>\-md12\, i10=>\-md13\, i9=>\-md14\, i8=>\-md15\, i7=>\-md16\);
  trap_1e30 : ic_93s48 port map(i6    => \-md29\, i5 => \-md30\, i4=>\-md31\, i3=>mdparl, i2=>mdparm, i1=>gnd, i0=>gnd, po=>mdparodd, pe=>mdpareven, i11=>\-md24\, i10=>\-md25\, i9=>\-md26\, i8=>\-md27\, i7=>\-md28\);
  trap_3e30 : ic_74s20 port map(g1a   => mdparerr, g1b => mdhaspar, g1c => \use.md\, g1d => \-wait\, g1y_n=>\-parerr\, g2a=>'0', g2b=>'0', g2c=>'0', g2d=>'0');
  trap_3f18 : ic_74s02 port map(g2q_n => \-trap\, g2a => internal17, g2b => \boot.trap\, g3b=>\-trapenb\, g3a=>\-parerr\, g3q_n=>internal17, g4b=>trapenb, g4a=>\-parerr\, g4q_n=>\-memparok\, g1a=>'0', g1b=>'0');
  trap_3f19 : ic_74s04 port map(g1a   => \-trap\, g1q_n => trapb, g2a => \-trap\, g2q_n=>trapa, g3a=>\-memparok\, g3q_n=>memparok, g4q=>\-trapenb\, g4a=>trapenb, g5a=>'0', g6a=>'0');

  spy0_1f01 : ic_74s138 port map(a => eadr0, b => eadr1, c => eadr2, g2a => \-dbread\, g2b => eadr3, g1 => hi1, y7 => \-spy.obh\, y6=>\-spy.obl\, y5=>\-spy.pc\, y4=>\-spy.opc\, y3=>nc3, y2=>\-spy.irh\, y1=>\-spy.irm\, y0=>\-spy.irl\);
  spy0_1f02 : ic_74s138 port map(a => eadr0, b => eadr1, c => eadr2, g2a => \-dbread\, g2b => gnd, g1 => eadr3, y7 => \-spy.sth\, y6=>\-spy.stl\, y5=>\-spy.ah\, y4=>\-spy.al\, y3=>\-spy.mh\, y2=>\-spy.ml\, y1=>\-spy.flag2\, y0=>\-spy.flag1\);
  spy0_1f03 : ic_74s138 port map(a => eadr0, b => eadr1, c => eadr2, g2a => \-dbwrite\, g2b => gnd, g1 => hi1, y7 => nc1, y6 => nc2, y5 => \-ldmode\, y4=>\-ldopc\, y3=>\-ldclk\, y2=>\-lddbirh\, y1=>\-lddbirm\, y0=>\-lddbirl\);

  spy1_2c17 : ic_74ls244 port map(aenb_n => \-spy.obl\, ain0 => ob7, bout3 => spy0, ain1 => ob6, bout2 => spy1, ain2 => ob5, bout1 => spy2, ain3 => ob4, bout0 => spy3, bin0 => ob3, aout3 => spy4, bin1 => ob2, aout2 => spy5, bin2 => ob1, aout1 => spy6, bin3 => ob0, aout0 => spy7, benb_n => \-spy.obl\);
  spy1_2c18 : ic_74ls244 port map(aenb_n => \-spy.obl\, ain0 => ob15, bout3 => spy8, ain1 => ob14, bout2 => spy9, ain2 => ob13, bout1 => spy10, ain3 => ob12, bout0 => spy11, bin0 => ob11, aout3 => spy12, bin1 => ob10, aout2 => spy13, bin2 => ob9, aout1 => spy14, bin3 => ob8, aout0 => spy15, benb_n => \-spy.obl\);
  spy1_3c23 : ic_74ls244 port map(aenb_n => \-spy.obh\, ain0 => ob23, bout3 => spy0, ain1 => ob22, bout2 => spy1, ain2 => ob21, bout1 => spy2, ain3 => ob20, bout0 => spy3, bin0 => ob19, aout3 => spy4, bin1 => ob18, aout2 => spy5, bin2 => ob17, aout1 => spy6, bin3 => ob16, aout0 => spy7, benb_n => \-spy.obh\);
  spy1_3c24 : ic_74ls244 port map(aenb_n => \-spy.obh\, ain0 => ob31, bout3 => spy8, ain1 => ob30, bout2 => spy9, ain2 => ob29, bout1 => spy10, ain3 => ob28, bout0 => spy11, bin0 => ob27, aout3 => spy12, bin1 => ob26, aout2 => spy13, bin2 => ob25, aout1 => spy14, bin3 => ob24, aout0 => spy15, benb_n => \-spy.obh\);
  spy1_3e01 : ic_74ls244 port map(aenb_n => \-spy.irl\, ain0 => ir7, bout3 => spy0, ain1 => ir6, bout2 => spy1, ain2 => ir5, bout1 => spy2, ain3 => ir4, bout0 => spy3, bin0 => ir3, aout3 => spy4, bin1 => ir2, aout2 => spy5, bin2 => ir1, aout1 => spy6, bin3 => ir0, aout0 => spy7, benb_n => \-spy.irl\);
  spy1_3e03 : ic_74ls244 port map(aenb_n => \-spy.irl\, ain0 => ir15, bout3 => spy8, ain1 => ir14, bout2 => spy9, ain2 => ir13, bout1 => spy10, ain3 => ir12, bout0 => spy11, bin0 => ir11, aout3 => spy12, bin1 => ir10, aout2 => spy13, bin2 => ir9, aout1 => spy14, bin3 => ir8, aout0 => spy15, benb_n => \-spy.irl\);
  spy1_3e06 : ic_74ls244 port map(aenb_n => \-spy.irh\, ain0 => ir47, bout3 => spy8, ain1 => ir46, bout2 => spy9, ain2 => ir45, bout1 => spy10, ain3 => ir44, bout0 => spy11, bin0 => ir43, aout3 => spy12, bin1 => ir42, aout2 => spy13, bin2 => ir41, aout1 => spy14, bin3 => ir40, aout0 => spy15, benb_n => \-spy.irh\);
  spy1_3f21 : ic_74ls244 port map(aenb_n => \-spy.irh\, ain0 => ir39, bout3 => spy0, ain1 => ir38, bout2 => spy1, ain2 => ir37, bout1 => spy2, ain3 => ir36, bout0 => spy3, bin0 => ir35, aout3 => spy4, bin1 => ir34, aout2 => spy5, bin2 => ir33, aout1 => spy6, bin3 => ir32, aout0 => spy7, benb_n => \-spy.irh\);
  spy1_3f23 : ic_74ls244 port map(aenb_n => \-spy.irm\, ain0 => ir31, bout3 => spy8, ain1 => ir30, bout2 => spy9, ain2 => ir29, bout1 => spy10, ain3 => ir28, bout0 => spy11, bin0 => ir27, aout3 => spy12, bin1 => ir26, aout2 => spy13, bin2 => ir25, aout1 => spy14, bin3 => ir24, aout0 => spy15, benb_n => \-spy.irm\);
  spy1_3f25 : ic_74ls244 port map(aenb_n => \-spy.irm\, ain0 => ir23, bout3 => spy0, ain1 => ir22, bout2 => spy1, ain2 => ir21, bout1 => spy2, ain3 => ir20, bout0 => spy3, bin0 => ir19, aout3 => spy4, bin1 => ir18, aout2 => spy5, bin2 => ir17, aout1 => spy6, bin3 => ir16, aout0 => spy7, benb_n => \-spy.irm\);

  spy2_1f11 : ic_74ls244 port map(aenb_n => \-spy.al\, ain0 => aa15, bout3 => spy8, ain1 => aa14, bout2 => spy9, ain2 => aa13, bout1 => spy10, ain3 => aa12, bout0 => spy11, bin0 => aa11, aout3 => spy12, bin1 => aa10, aout2 => spy13, bin2 => aa9, aout1 => spy14, bin3 => aa8, aout0 => spy15, benb_n => \-spy.al\);
  spy2_1f13 : ic_74ls244 port map(aenb_n => \-spy.al\, ain0 => aa7, bout3 => spy0, ain1 => aa6, bout2 => spy1, ain2 => aa5, bout1 => spy2, ain3 => aa4, bout0 => spy3, bin0 => aa3, aout3 => spy4, bin1 => aa2, aout2 => spy5, bin2 => aa1, aout1 => spy6, bin3 => aa0, aout0 => spy7, benb_n => \-spy.al\);
  spy2_3a26 : ic_74ls244 port map(aenb_n => \-spy.ah\, ain0 => a31a, bout3 => spy8, ain1 => a30, bout2 => spy9, ain2 => a29, bout1 => spy10, ain3 => a28, bout0 => spy11, bin0 => a27, aout3 => spy12, bin1 => a26, aout2 => spy13, bin2 => a25, aout1 => spy14, bin3 => a24, aout0 => spy15, benb_n => \-spy.ah\);
  spy2_3a27 : ic_74ls244 port map(aenb_n => \-spy.ah\, ain0 => a23, bout3 => spy0, ain1 => a22, bout2 => spy1, ain2 => a21, bout1 => spy2, ain3 => a20, bout0 => spy3, bin0 => a19, aout3 => spy4, bin1 => a18, aout2 => spy5, bin2 => a17, aout1 => spy6, bin3 => a16, aout0 => spy7, benb_n => \-spy.ah\);
  spy2_3e16 : ic_74ls244 port map(aenb_n => \-spy.flag2\, ain0 => nc149, bout3 => spy0, ain1 => nc150, bout2 => spy1, ain2 => ir48, bout1 => spy2, ain3 => nop, bout0 => spy3, bin0 => \-vmaok\, aout3=>spy4, bin1=>jcond, aout2=>spy5, bin2=>pcs1, aout1=>spy6, bin3=>pcs0, aout0=>spy7, benb_n=>\-spy.flag2\);
  spy2_3f15 : ic_74ls244 port map(aenb_n => \-spy.flag2\, ain0 => nc151, bout3 => spy8, ain1 => nc152, bout2 => spy9, ain2 => wmapd, bout1 => spy10, ain3 => destspcd, bout0 => spy11, bin0 => iwrited, aout3 => spy12, bin1 => imodd, aout2 => spy13, bin2 => pdlwrited, aout1 => spy14, bin3 => spushd, aout0 => spy15, benb_n => \-spy.flag2\);
  spy2_4a13 : ic_74ls244 port map(aenb_n => \-spy.ml\, ain0 => m15, bout3 => spy8, ain1 => m14, bout2 => spy9, ain2 => m13, bout1 => spy10, ain3 => m12, bout0 => spy11, bin0 => m11, aout3 => spy12, bin1 => m10, aout2 => spy13, bin2 => m9, aout1 => spy14, bin3 => m8, aout0 => spy15, benb_n => \-spy.ml\);
  spy2_4a15 : ic_74ls244 port map(aenb_n => \-spy.ml\, ain0 => m7, bout3 => spy0, ain1 => m6, bout2 => spy1, ain2 => m5, bout1 => spy2, ain3 => m4, bout0 => spy3, bin0 => m3, aout3 => spy4, bin1 => m2, aout2 => spy5, bin2 => m1, aout1 => spy6, bin3 => m0, aout0 => spy7, benb_n => \-spy.ml\);
  spy2_4b13 : ic_74ls244 port map(aenb_n => \-spy.mh\, ain0 => m23, bout3 => spy0, ain1 => m22, bout2 => spy1, ain2 => m21, bout1 => spy2, ain3 => m20, bout0 => spy3, bin0 => m19, aout3 => spy4, bin1 => m18, aout2 => spy5, bin2 => m17, aout1 => spy6, bin3 => m16, aout0 => spy7, benb_n => \-spy.mh\);
  spy2_4b17 : ic_74ls244 port map(aenb_n => \-spy.mh\, ain0 => m31, bout3 => spy8, ain1 => m30, bout2 => spy9, ain2 => m29, bout1 => spy10, ain3 => m28, bout0 => spy11, bin0 => m27, aout3 => spy12, bin1 => m26, aout2 => spy13, bin2 => m25, aout1 => spy14, bin3 => m24, aout0 => spy15, benb_n => \-spy.mh\);

  spy4_1a12 : ic_74ls244 port map(aenb_n => \-spy.flag1\, ain0 => \-wait\, bout3=>spy8, ain1=>\-v1pe\, bout2=>spy9, ain2=>\-v0pe\, bout1=>spy10, ain3=>promdisable, bout0=>spy11, bin0=>\-stathalt\, aout3=>spy12, bin1=>err, aout2=>spy13, bin2=>ssdone, aout1=>spy14, bin3=>srun, aout0=>spy15, benb_n=>\-spy.flag1\);
  spy4_1a13 : ic_74s240 port map(aenb_n  => \-spy.flag1\, ain0 => \-higherr\, bout3=>spy0, ain1=>\-mempe\, bout2=>spy1, ain2=>\-ipe\, bout1=>spy2, ain3=>\-dpe\, bout0=>spy3, bin0=>\-spe\, aout3=>spy4, bin1=>\-pdlpe\, aout2=>spy5, bin2=>\-mpe\, aout1=>spy6, bin3=>\-ape\, aout0=>spy7, benb_n=>\-spy.flag1\);
  spy4_1d06 : ic_74ls244 port map(aenb_n => \-spy.pc\, ain0 => gnd, bout3 => spy8, ain1 => gnd, bout2 => spy9, ain2 => pc13, bout1 => spy10, ain3 => pc12, bout0 => spy11, bin0 => pc11, aout3 => spy12, bin1 => pc10, aout2 => spy13, bin2 => pc9, aout1 => spy14, bin3 => pc8, aout0 => spy15, benb_n => \-spy.pc\);
  spy4_1d07 : ic_74ls244 port map(aenb_n => \-spy.pc\, ain0 => pc7, bout3 => spy0, ain1 => pc6, bout2 => spy1, ain2 => pc5, bout1 => spy2, ain3 => pc4, bout0 => spy3, bin0 => pc3, aout3 => spy4, bin1 => pc2, aout2 => spy5, bin2 => pc1, aout1 => spy6, bin3 => pc0, aout0 => spy7, benb_n => \-spy.pc\);
  spy4_1e06 : ic_74ls244 port map(aenb_n => \-spy.opc\, ain0 => gnd, bout3 => spy8, ain1 => gnd, bout2 => spy9, ain2 => opc13, bout1 => spy10, ain3 => opc12, bout0 => spy11, bin0 => opc11, aout3 => spy12, bin1 => opc10, aout2 => spy13, bin2 => opc9, aout1 => spy14, bin3 => opc8, aout0 => spy15, benb_n => \-spy.opc\);
  spy4_1e07 : ic_74ls244 port map(aenb_n => \-spy.opc\, ain0 => opc7, bout3 => spy0, ain1 => opc6, bout2 => spy1, ain2 => opc5, bout1 => spy2, ain3 => opc4, bout0 => spy3, bin0 => opc3, aout3 => spy4, bin1 => opc2, aout2 => spy5, bin2 => opc1, aout1 => spy6, bin3 => opc0, aout0 => spy7, benb_n => \-spy.opc\);

  opcd_1d18 : ic_74s04 port map(g2a     => \-srcdc\, g2q_n => internal20, g3a => \-srcopc\, g3q_n=>internal21, g1a=>'0', g4a=>'0', g5a=>'0', g6a=>'0');
  opcd_1e01 : ic_74s241 port map(aenb_n => \-opcdrive\, ain0 => opc7, bout3 => mf4, ain1 => opc6, bout2 => mf5, ain2 => opc5, bout1 => mf6, ain3 => opc4, bout0 => mf7, bin0 => dc7, aout3 => mf4, bin1 => dc6, aout2 => mf5, bin2 => dc5, aout1 => mf6, bin3 => dc4, aout0 => mf7, benb => dcdrive);
  opcd_1e03 : ic_74s241 port map(aenb_n => \-opcdrive\, ain0 => opc3, bout3 => mf0, ain1 => opc2, bout2 => mf1, ain2 => opc1, bout1 => mf2, ain3 => opc0, bout0 => mf3, bin0 => dc3, aout3 => mf0, bin1 => dc2, aout2 => mf1, bin2 => dc1, aout1 => mf2, bin3 => dc0, aout0 => mf3, benb => dcdrive);
  opcd_1e06 : ic_74s00 port map(g3q_n   => \-opcdrive\, g3b => internal21, g3a => tse1b, g4q_n => \-zero16.drive\, g4a=>tse1b, g4b=>zero16, g1b=>'0', g1a=>'0', g2b=>'0', g2a=>'0');
  opcd_1e07 : ic_74s08 port map(g1b     => tse1b, g1a => internal20, g1q => dcdrive, g2b => zero16, g2a => tse1b, g2q => \zero16.drive\, g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  opcd_1e16 : ic_74s11 port map(g1a     => \-srcopc\, g1b => zero16, g1y_n => \zero12.drive\, g1c=>tse1b, g2a=>'0', g2b=>'0', g2c=>'0', g3a=>'0', g3b=>'0', g3c=>'0');
  opcd_1f01 : ic_74s241 port map(aenb_n => \-zero16.drive\, ain0 => gnd, bout3 => mf24, ain1 => gnd, bout2 => mf25, ain2 => gnd, bout1 => mf26, ain3 => gnd, bout0 => mf27, bin0 => gnd, aout3 => mf28, bin1 => gnd, aout2 => mf29, bin2 => gnd, aout1 => mf30, bin3 => gnd, aout0 => mf31, benb => \zero16.drive\);
  opcd_1f02 : ic_74s241 port map(aenb_n => \-zero16.drive\, ain0 => gnd, bout3 => mf16, ain1 => gnd, bout2 => mf17, ain2 => gnd, bout1 => mf18, ain3 => gnd, bout0 => mf19, bin0 => gnd, aout3 => mf20, bin1 => gnd, aout2 => mf21, bin2 => gnd, aout1 => mf22, bin3 => gnd, aout0 => mf23, benb => \zero16.drive\);
  opcd_1f03 : ic_74s241 port map(aenb_n => \-opcdrive\, ain0 => gnd, bout3 => mf12, ain1 => gnd, bout2 => mf13, ain2 => opc13, bout1 => mf14, ain3 => opc12, bout0 => mf15, bin0 => gnd, aout3 => mf12, bin1 => gnd, aout2 => mf13, bin2 => gnd, aout1 => mf14, bin3 => gnd, aout0 => mf15, benb => \zero12.drive\);
  opcd_1f04 : ic_74s241 port map(aenb_n => \-opcdrive\, ain0 => opc11, bout3 => mf8, ain1 => opc10, bout2 => mf9, ain2 => opc9, bout1 => mf10, ain3 => opc8, bout0 => mf11, bin0 => gnd, aout3 => mf8, bin1 => gnd, aout2 => mf9, bin2 => dc9, aout1 => mf10, bin3 => dc8, aout0 => mf11, benb => dcdrive);
  opcd_3e30 : ic_74s20 port map(g2y_n   => zero16, g2a => \-srcopc\, g2b => \-srcpdlidx\, g2c=>\-srcpdlptr\, g2d=>\-srcdc\, g1a=>'0', g1b=>'0', g1c=>'0', g1d=>'0');

  mo0_2a24 : ic_74s151 port map(i3 => alu15, i2 => alu15, i1 => r15, i0 => a15, q => ob15, q_n => nc290, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk15, i7 => alu14, i6 => alu14, i5 => alu16, i4 => alu16);
  mo0_2a25 : ic_74s151 port map(i3 => alu14, i2 => alu14, i1 => r14, i0 => a14, q => ob14, q_n => nc289, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk14, i7 => alu13, i6 => alu13, i5 => alu15, i4 => alu15);
  mo0_2a29 : ic_74s151 port map(i3 => alu13, i2 => alu13, i1 => r13, i0 => a13, q => ob13, q_n => nc288, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk13, i7 => alu12, i6 => alu12, i5 => alu14, i4 => alu14);
  mo0_2a30 : ic_74s151 port map(i3 => alu12, i2 => alu12, i1 => r12, i0 => a12, q => ob12, q_n => nc287, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk12, i7 => alu11, i6 => alu11, i5 => alu13, i4 => alu13);
  mo0_2b24 : ic_74s151 port map(i3 => alu7, i2 => alu7, i1 => r7, i0 => a7, q => ob7, q_n => nc282, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk7, i7 => alu6, i6 => alu6, i5 => alu8, i4 => alu8);
  mo0_2b25 : ic_74s151 port map(i3 => alu6, i2 => alu6, i1 => r6, i0 => a6, q => ob6, q_n => nc281, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk6, i7 => alu5, i6 => alu5, i5 => alu7, i4 => alu7);
  mo0_2b29 : ic_74s151 port map(i3 => alu5, i2 => alu5, i1 => r5, i0 => a5, q => ob5, q_n => nc280, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk5, i7 => alu4, i6 => alu4, i5 => alu6, i4 => alu6);
  mo0_2b30 : ic_74s151 port map(i3 => alu4, i2 => alu4, i1 => r4, i0 => a4, q => ob4, q_n => nc279, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk4, i7 => alu3, i6 => alu3, i5 => alu5, i4 => alu5);
  mo0_2c19 : ic_74s151 port map(i3 => alu11, i2 => alu11, i1 => r11, i0 => a11, q => ob11, q_n => nc286, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk11, i7 => alu10, i6 => alu10, i5 => alu12, i4 => alu12);
  mo0_2c24 : ic_74s151 port map(i3 => alu10, i2 => alu10, i1 => r10, i0 => a10, q => ob10, q_n => nc285, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk10, i7 => alu9, i6 => alu9, i5 => alu11, i4 => alu11);
  mo0_2c29 : ic_74s151 port map(i3 => alu3, i2 => alu3, i1 => r3, i0 => a3, q => ob3, q_n => nc278, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk3, i7 => alu2, i6 => alu2, i5 => alu4, i4 => alu4);
  mo0_2c30 : ic_74s151 port map(i3 => alu2, i2 => alu2, i1 => r2, i0 => a2, q => ob2, q_n => nc277, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk2, i7 => alu1, i6 => alu1, i5 => alu3, i4 => alu3);
  mo0_2d23 : ic_74s151 port map(i3 => alu9, i2 => alu9, i1 => r9, i0 => a9, q => ob9, q_n => nc284, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk9, i7 => alu8, i6 => alu8, i5 => alu10, i4 => alu10);
  mo0_2d24 : ic_74s151 port map(i3 => alu8, i2 => alu8, i1 => r8, i0 => a8, q => ob8, q_n => nc283, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk8, i7 => alu7, i6 => alu7, i5 => alu9, i4 => alu9);
  mo0_2d28 : ic_74s151 port map(i3 => alu1, i2 => alu1, i1 => r1, i0 => a1, q => ob1, q_n => nc276, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk1, i7 => alu0, i6 => alu0, i5 => alu2, i4 => alu2);
  mo0_2d29 : ic_74s151 port map(i3 => alu0, i2 => alu0, i1 => r0, i0 => a0, q => ob0, q_n => nc275, ce_n => gnd, sel2 => osel1b, sel1 => osel0b, sel0 => msk0, i7 => q31, i6 => q31, i5 => alu1, i4 => alu1);

  mo1_2a09 : ic_74s151 port map(i3 => alu31, i2 => alu31, i1 => r31, i0 => a31b, q => ob31, q_n => nc274, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk31, i7 => alu30, i6 => alu30, i5 => alu32, i4 => alu32);
  mo1_2a10 : ic_74s151 port map(i3 => alu30, i2 => alu30, i1 => r30, i0 => a30, q => ob30, q_n => nc273, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk30, i7 => alu29, i6 => alu29, i5 => alu31, i4 => alu31);
  mo1_2a14 : ic_74s151 port map(i3 => alu29, i2 => alu29, i1 => r29, i0 => a29, q => ob29, q_n => nc272, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk29, i7 => alu28, i6 => alu28, i5 => alu30, i4 => alu30);
  mo1_2a15 : ic_74s151 port map(i3 => alu28, i2 => alu28, i1 => r28, i0 => a28, q => ob28, q_n => nc271, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk28, i7 => alu27, i6 => alu27, i5 => alu29, i4 => alu29);
  mo1_2b09 : ic_74s151 port map(i3 => alu23, i2 => alu23, i1 => r23, i0 => a23, q => ob23, q_n => nc266, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk23, i7 => alu22, i6 => alu22, i5 => alu24, i4 => alu24);
  mo1_2b10 : ic_74s151 port map(i3 => alu22, i2 => alu22, i1 => r22, i0 => a22, q => ob22, q_n => nc265, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk22, i7 => alu21, i6 => alu21, i5 => alu23, i4 => alu23);
  mo1_2b14 : ic_74s151 port map(i3 => alu21, i2 => alu21, i1 => r21, i0 => a21, q => ob21, q_n => nc264, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk21, i7 => alu20, i6 => alu20, i5 => alu22, i4 => alu22);
  mo1_2b15 : ic_74s151 port map(i3 => alu20, i2 => alu20, i1 => r20, i0 => a20, q => ob20, q_n => nc263, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk20, i7 => alu19, i6 => alu19, i5 => alu21, i4 => alu21);
  mo1_2c09 : ic_74s151 port map(i3 => alu27, i2 => alu27, i1 => r27, i0 => a27, q => ob27, q_n => nc270, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk27, i7 => alu26, i6 => alu26, i5 => alu28, i4 => alu28);
  mo1_2c14 : ic_74s151 port map(i3 => alu24, i2 => alu24, i1 => r24, i0 => a24, q => ob24, q_n => nc267, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk24, i7 => alu23, i6 => alu23, i5 => alu25, i4 => alu25);
  mo1_2d04 : ic_74s151 port map(i3 => alu26, i2 => alu26, i1 => r26, i0 => a26, q => ob26, q_n => nc269, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk26, i7 => alu25, i6 => alu25, i5 => alu27, i4 => alu27);
  mo1_2d09 : ic_74s151 port map(i3 => alu25, i2 => alu25, i1 => r25, i0 => a25, q => ob25, q_n => nc268, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk25, i7 => alu24, i6 => alu24, i5 => alu26, i4 => alu26);
  mo1_2d13 : ic_74s151 port map(i3 => alu19, i2 => alu19, i1 => r19, i0 => a19, q => ob19, q_n => nc262, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk19, i7 => alu18, i6 => alu18, i5 => alu20, i4 => alu20);
  mo1_2d14 : ic_74s151 port map(i3 => alu18, i2 => alu18, i1 => r18, i0 => a18, q => ob18, q_n => nc261, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk18, i7 => alu17, i6 => alu17, i5 => alu19, i4 => alu19);
  mo1_2d18 : ic_74s151 port map(i3 => alu17, i2 => alu17, i1 => r17, i0 => a17, q => ob17, q_n => nc260, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk17, i7 => alu16, i6 => alu16, i5 => alu18, i4 => alu18);
  mo1_2d19 : ic_74s151 port map(i3 => alu16, i2 => alu16, i1 => r16, i0 => a16, q => ob16, q_n => nc259, ce_n => gnd, sel2 => osel1a, sel1 => osel0a, sel0 => msk16, i7 => alu15, i6 => alu15, i5 => alu17, i4 => alu17);

  bcterm_1b15 : ic_sip220_330_8 port map(r2 => mem0, r3 => mem1, r4 => mem2, r5 => mem3, r6 => mem4, r7 => mem5);
  bcterm_1b20 : ic_sip220_330_8 port map(r2 => mem12, r3 => mem13, r4 => mem14, r5 => mem15, r6 => mem16, r7 => mem17);
  bcterm_1b25 : ic_sip220_330_8 port map(r2 => mem24, r3 => mem25, r4 => mem26, r5 => mem27, r6 => mem28, r7 => mem29);
  bcterm_2c25 : ic_sip330_470_8 port map(r2 => \-memgrant\, r3 => int, r4 => \-loadmd\, r5=>\-ignpar\, r6=>\-memack\, r7=>nc431);

  ipar_3e02 : ic_93s48 port map(i6  => ir41, i5 => ir42, i4 => ir43, i3 => ir44, i2 => ir45, i1 => ir46, i0 => ir47, po => ipar3, pe => nc381, i11 => ir36, i10 => ir37, i9 => ir38, i8 => ir39, i7 => ir40);
  ipar_3e04 : ic_93s48 port map(i6  => ir5, i5 => ir6, i4 => ir7, i3 => ir8, i2 => ir9, i1 => ir10, i0 => ir11, po => ipar0, pe => nc384, i11 => ir0, i10 => ir1, i9 => ir2, i8 => ir3, i7 => ir4);
  ipar_3e21 : ic_93s48 port map(i6  => ir29, i5 => ir30, i4 => ir31, i3 => ir32, i2 => ir33, i1 => ir34, i0 => ir35, po => ipar2, pe => nc382, i11 => ir24, i10 => ir25, i9 => ir26, i8 => ir27, i7 => ir28);
  ipar_3f22 : ic_93s48 port map(i6  => gnd, i5 => gnd, i4 => gnd, i3 => gnd, i2 => gnd, i1 => gnd, i0 => gnd, po => iparity, pe => nc380, i11 => ipar0, i10 => ipar1, i9 => ipar2, i8 => ipar3, i7 => ir48);
  ipar_3f24 : ic_93s48 port map(i6  => ir17, i5 => ir18, i4 => ir19, i3 => ir20, i2 => ir21, i1 => ir22, i0 => ir23, po => ipar1, pe => nc383, i11 => ir12, i10 => ir13, i9 => ir14, i8 => ir15, i7 => ir16);
  ipar_4e03 : ic_74s32 port map(g2a => imodd, g2b => iparity, g2y => iparok, g1a => '0', g1b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');

  --------------------------------------------------------------------------------

  -- Poor substitute for the 5 octal display that was on the lower
  -- left-hand corner of the front door on the CADR.  See the PCTL
  -- prints.
  process (cyclecompleted)
  begin
    pc <= pc0 & pc1 & pc2 & pc3 & pc4 & pc5 & pc6 & pc7 & pc8 & pc9 & pc10 & pc12 & pc13;

    report "PC: " & to_hstring(pc);
    if tilt1 then report "TILT1"; end if;
    if tilt0 then report "TILT0"; end if;
    if dpe then report "DPE"; end if;
    if ipe then report "IPE"; end if;
    if promenable then report "PROMENABLE"; end if;
  end process;

  process
  begin
    wait for 0.1 ns;
  end process;

end;
