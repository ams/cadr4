library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_olord1 is
  port (
    \-clock_reset_a\ : in  std_logic;
    speed1a          : out std_logic;
    sspeed1          : out std_logic;
    speedclk         : out std_logic;
    sspeed0          : out std_logic;
    speed0a          : out std_logic;
    speed1           : out std_logic;
    speed0           : out std_logic;
    \-reset\         : in  std_logic;
    spy0             : in  std_logic;
    spy1             : in  std_logic;
    spy2             : in  std_logic;
    errstop          : out std_logic;
    \-ldmode\        : in  std_logic;
    stathenb         : out std_logic;
    spy3             : in  std_logic;
    trapenb          : out std_logic;
    spy4             : in  std_logic;
    spy5             : in  std_logic;
    promdisable      : out std_logic;
    \-opcinh\        : out std_logic;
    opcinh           : out std_logic;
    \-ldopc\         : in  std_logic;
    opcclk           : out std_logic;
    \-opcclk\        : out std_logic;
    \-lpc.hold\      : out std_logic;
    \lpc.hold\       : out std_logic;
    ldstat           : out std_logic;
    \-ldstat\        : out std_logic;
    \-idebug\        : out std_logic;
    idebug           : out std_logic;
    \-ldclk\         : in  std_logic;
    nop11            : out std_logic;
    \-nop11\         : out std_logic;
    \-step\          : out std_logic;
    step             : out std_logic;
    promdisabled     : out std_logic;
    sstep            : out std_logic;
    ssdone           : out std_logic;
    mclk5a           : in  std_logic;
    srun             : out std_logic;
    run              : out std_logic;
    \-boot\          : in  std_logic;
    \-run\           : out std_logic;
    \-ssdone\        : out std_logic;
    \-errhalt\       : in  std_logic;
    \-wait\          : in  std_logic;
    \-stathalt\      : out std_logic;
    machrun          : out std_logic;
    \stat.ovf\       : out std_logic;
    \-stc32\         : in  std_logic;
    \-tpr60\         : in  std_logic;
    gnd              : in  std_logic;
    statstop         : in  std_logic;
    \-machruna\      : out std_logic;
    \-machrun\       : out std_logic);
end;

architecture ttl of cadr4_olord1 is
  signal nc84 : std_logic;
  signal nc85 : std_logic;
  signal nc86 : std_logic;
  signal nc87 : std_logic;
  signal nc88 : std_logic;
  signal nc89 : std_logic;
  signal nc90 : std_logic;
  signal nc91 : std_logic;
  signal nc92 : std_logic;
  signal nc93 : std_logic;
begin
  olord1_1a01 : sn74s174 port map(clr_n => \-clock_reset_a\, q1 => nc84, d1 => nc85, d2 => nc86, q2 => nc87, d3 => speed1a, q3 => sspeed1, clk => speedclk, q4 => sspeed0, d4 => speed0a, q5 => speed1a, d5 => speed1, d6 => speed0, q6 => speed0a);
  olord1_1a04 : sn74s174 port map(clr_n => \-reset\, q1 => speed0, d1 => spy0, d2 => spy1, q2 => speed1, d3 => spy2, q3 => errstop, clk => \-ldmode\, q4 => stathenb, d4 => spy3, q5 => trapenb, d5 => spy4, d6 => spy5, q6 => promdisable);
  olord1_1a08 : sn74s175 port map(clr_n => \-reset\, q0 => nc92, q0_n => nc93, d0 => spy3, d1 => spy2, q1_n => \-opcinh\, q1 => opcinh, clk => \-ldopc\, q2 => opcclk, q2_n => \-opcclk\, d2 => spy1, d3 => spy0, q3_n => \-lpc.hold\, q3 => \lpc.hold\);
  olord1_1a09 : sn74s175 port map(clr_n => \-reset\, q0 => ldstat, q0_n => \-ldstat\, d0 => spy4, d1 => spy3, q1_n => \-idebug\, q1 => idebug, clk => \-ldclk\, q2 => nop11, q2_n => \-nop11\, d2 => spy2, d3 => spy1, q3_n => \-step\, q3 => step);
  olord1_1a10 : sn74s174 port map(clr_n => \-clock_reset_a\, q1 => promdisabled, d1 => promdisable, d2 => sstep, q2 => ssdone, d3 => step, q3 => sstep, clk => mclk5a, q4 => srun, d4 => run, q5 => nc88, d5 => nc89, d6 => nc90, q6 => nc91);
  olord1_1a14 : sn74s74 port map(g1r_n  => \-clock_reset_a\, g1d => spy0, g1clk => \-ldclk\, g1s_n => \-boot\, g1q => run, g1q_n => \-run\, g2s_n => '0', g2clk => '0', g2d => '0', g2r_n => '0');
  olord1_1a15 : dm9s42_1 port map(g1a1  => sstep, g1b1 => \-ssdone\, g2a1 => srun, g2b1 => \-errhalt\, g2c1 => \-wait\, g2d1 => \-stathalt\, out1 => machrun, g1a2 => '0', g1b2 => '0', g2a2 => '0', g2b2 => '0', g2c2 => '0', g2d2 => '0');
  olord1_1b10 : sn74s04 port map(g2a    => ssdone, g2q_n => \-ssdone\, g5q_n => \stat.ovf\, g5a => \-stc32\, g1a => '0', g3a => '0', g4a => '0', g6a => '0');
  olord1_1c01 : sn7428 port map(g3a     => \-tpr60\, g3b => gnd, g3q_n => speedclk, g1a => '0', g1b => '0', g2a => '0', g4a => '0', g4b => '0', g2b => '0');
  olord1_1c09 : sn74s00 port map(g3q_n  => \-stathalt\, g3b => stathenb, g3a => statstop, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  olord1_1c10 : sn74s02 port map(g1q_n  => \-machruna\, g1a => gnd, g1b => machrun, g2a => '0', g2b => '0', g3b => '0', g3a => '0', g4b => '0', g4a => '0');
  olord1_1f10 : sn74s04 port map(g4q_n  => \-machrun\, g4a => machrun, g1a => '0', g2a => '0', g3a => '0', g5a => '0', g6a => '0');
end architecture;
