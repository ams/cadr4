library ieee;
use ieee.std_logic_1164.all;

entity cadr_mlatch is
  port (
    \-mpassl\       : in     std_logic;
    \-mpassm\       : in     std_logic;
    clk4a           : in     std_logic;
    l0              : in     std_logic;
    l1              : in     std_logic;
    l10             : in     std_logic;
    l11             : in     std_logic;
    l12             : in     std_logic;
    l13             : in     std_logic;
    l14             : in     std_logic;
    l15             : in     std_logic;
    l16             : in     std_logic;
    l17             : in     std_logic;
    l18             : in     std_logic;
    l19             : in     std_logic;
    l2              : in     std_logic;
    l20             : in     std_logic;
    l21             : in     std_logic;
    l22             : in     std_logic;
    l23             : in     std_logic;
    l24             : in     std_logic;
    l25             : in     std_logic;
    l26             : in     std_logic;
    l27             : in     std_logic;
    l28             : in     std_logic;
    l29             : in     std_logic;
    l3              : in     std_logic;
    l30             : in     std_logic;
    l31             : in     std_logic;
    l4              : in     std_logic;
    l5              : in     std_logic;
    l6              : in     std_logic;
    l7              : in     std_logic;
    l8              : in     std_logic;
    l9              : in     std_logic;
    mmem0           : in     std_logic;
    mmem1           : in     std_logic;
    mmem10          : in     std_logic;
    mmem11          : in     std_logic;
    mmem12          : in     std_logic;
    mmem13          : in     std_logic;
    mmem14          : in     std_logic;
    mmem15          : in     std_logic;
    mmem16          : in     std_logic;
    mmem17          : in     std_logic;
    mmem18          : in     std_logic;
    mmem19          : in     std_logic;
    mmem2           : in     std_logic;
    mmem20          : in     std_logic;
    mmem21          : in     std_logic;
    mmem22          : in     std_logic;
    mmem23          : in     std_logic;
    mmem24          : in     std_logic;
    mmem25          : in     std_logic;
    mmem26          : in     std_logic;
    mmem27          : in     std_logic;
    mmem28          : in     std_logic;
    mmem29          : in     std_logic;
    mmem3           : in     std_logic;
    mmem30          : in     std_logic;
    mmem31          : in     std_logic;
    mmem4           : in     std_logic;
    mmem5           : in     std_logic;
    mmem6           : in     std_logic;
    mmem7           : in     std_logic;
    mmem8           : in     std_logic;
    mmem9           : in     std_logic;
    mmemparity      : in     std_logic;
    mpassl          : in     std_logic;
    m0              : out    std_logic;
    m1              : out    std_logic;
    m10             : out    std_logic;
    m11             : out    std_logic;
    m12             : out    std_logic;
    m13             : out    std_logic;
    m14             : out    std_logic;
    m15             : out    std_logic;
    m16             : out    std_logic;
    m17             : out    std_logic;
    m18             : out    std_logic;
    m19             : out    std_logic;
    m2              : out    std_logic;
    m20             : out    std_logic;
    m21             : out    std_logic;
    m22             : out    std_logic;
    m23             : out    std_logic;
    m24             : out    std_logic;
    m25             : out    std_logic;
    m26             : out    std_logic;
    m27             : out    std_logic;
    m28             : out    std_logic;
    m29             : out    std_logic;
    m3              : out    std_logic;
    m30             : out    std_logic;
    m31             : out    std_logic;
    m4              : out    std_logic;
    m5              : out    std_logic;
    m6              : out    std_logic;
    m7              : out    std_logic;
    m8              : out    std_logic;
    m9              : out    std_logic;
    mf0             : out    std_logic;
    mf1             : out    std_logic;
    mf10            : out    std_logic;
    mf11            : out    std_logic;
    mf12            : out    std_logic;
    mf13            : out    std_logic;
    mf14            : out    std_logic;
    mf15            : out    std_logic;
    mf16            : out    std_logic;
    mf17            : out    std_logic;
    mf18            : out    std_logic;
    mf19            : out    std_logic;
    mf2             : out    std_logic;
    mf20            : out    std_logic;
    mf21            : out    std_logic;
    mf22            : out    std_logic;
    mf23            : out    std_logic;
    mf24            : out    std_logic;
    mf25            : out    std_logic;
    mf26            : out    std_logic;
    mf27            : out    std_logic;
    mf28            : out    std_logic;
    mf29            : out    std_logic;
    mf3             : out    std_logic;
    mf30            : out    std_logic;
    mf31            : out    std_logic;
    mf4             : out    std_logic;
    mf5             : out    std_logic;
    mf6             : out    std_logic;
    mf7             : out    std_logic;
    mf8             : out    std_logic;
    mf9             : out    std_logic;
    mparity         : out    std_logic
  );
end entity;
