library ieee;
use ieee.std_logic_1164.all;

use work.cadr_book.all;
use work.helper.all;
use work.icmem_book.all;

entity cadr_tb is
end entity;

architecture structural of cadr_tb is
  signal a0: std_logic;
  signal a1: std_logic;
  signal a2: std_logic;
  signal a3: std_logic;
  signal a4: std_logic;
  signal a5: std_logic;
  signal a6: std_logic;
  signal a7: std_logic;
  signal a8: std_logic;
  signal a9: std_logic;
  signal a10: std_logic;
  signal a11: std_logic;
  signal a12: std_logic;
  signal a13: std_logic;
  signal a14: std_logic;
  signal a15: std_logic;
  signal a16: std_logic;
  signal a17: std_logic;
  signal a18: std_logic;
  signal a19: std_logic;
  signal a20: std_logic;
  signal a21: std_logic;
  signal a22: std_logic;
  signal a23: std_logic;
  signal a24: std_logic;
  signal a25: std_logic;
  signal a26: std_logic;
  signal a27: std_logic;
  signal a28: std_logic;
  signal a29: std_logic;
  signal a30: std_logic;
  signal \-a31\: std_logic;
  signal a31a: std_logic;
  signal a31b: std_logic;
  signal \a=m\: std_logic;
  signal aa0: std_logic;
  signal aa1: std_logic;
  signal aa2: std_logic;
  signal aa3: std_logic;
  signal aa4: std_logic;
  signal aa5: std_logic;
  signal aa6: std_logic;
  signal aa7: std_logic;
  signal aa8: std_logic;
  signal aa9: std_logic;
  signal aa10: std_logic;
  signal aa11: std_logic;
  signal aa12: std_logic;
  signal aa13: std_logic;
  signal aa14: std_logic;
  signal aa15: std_logic;
  signal aa16: std_logic;
  signal aa17: std_logic;
  signal \-aadr0a\: std_logic;
  signal \-aadr0b\: std_logic;
  signal \-aadr1a\: std_logic;
  signal \-aadr1b\: std_logic;
  signal \-aadr2a\: std_logic;
  signal \-aadr2b\: std_logic;
  signal \-aadr3a\: std_logic;
  signal \-aadr3b\: std_logic;
  signal \-aadr4a\: std_logic;
  signal \-aadr4b\: std_logic;
  signal \-aadr5a\: std_logic;
  signal \-aadr5b\: std_logic;
  signal \-aadr6a\: std_logic;
  signal \-aadr6b\: std_logic;
  signal \-aadr7a\: std_logic;
  signal \-aadr7b\: std_logic;
  signal \-aadr8a\: std_logic;
  signal \-aadr8b\: std_logic;
  signal \-aadr9a\: std_logic;
  signal \-aadr9b\: std_logic;
  signal \-adrpar\: std_logic;
  signal alu0: std_logic;
  signal alu1: std_logic;
  signal alu2: std_logic;
  signal alu3: std_logic;
  signal alu4: std_logic;
  signal alu5: std_logic;
  signal alu6: std_logic;
  signal alu7: std_logic;
  signal alu8: std_logic;
  signal alu9: std_logic;
  signal alu10: std_logic;
  signal alu11: std_logic;
  signal alu12: std_logic;
  signal alu13: std_logic;
  signal alu14: std_logic;
  signal alu15: std_logic;
  signal alu16: std_logic;
  signal alu17: std_logic;
  signal alu18: std_logic;
  signal alu19: std_logic;
  signal alu20: std_logic;
  signal alu21: std_logic;
  signal alu22: std_logic;
  signal alu23: std_logic;
  signal alu24: std_logic;
  signal alu25: std_logic;
  signal alu26: std_logic;
  signal alu27: std_logic;
  signal alu28: std_logic;
  signal alu29: std_logic;
  signal alu30: std_logic;
  signal alu31: std_logic;
  signal \-alu31\: std_logic;
  signal alu32: std_logic;
  signal \-alu32\: std_logic;
  signal aluadd: std_logic;
  signal \-aluf0\: std_logic;
  signal \-aluf1\: std_logic;
  signal \-aluf2\: std_logic;
  signal \-aluf3\: std_logic;
  signal aluf0a: std_logic;
  signal aluf0b: std_logic;
  signal aluf1a: std_logic;
  signal aluf1b: std_logic;
  signal aluf2a: std_logic;
  signal aluf2b: std_logic;
  signal aluf3a: std_logic;
  signal aluf3b: std_logic;
  signal alumode: std_logic;
  signal \-alumode\: std_logic;
  signal aluneg: std_logic;
  signal alusub: std_logic;
  signal amem0: std_logic;
  signal amem1: std_logic;
  signal amem2: std_logic;
  signal amem3: std_logic;
  signal amem4: std_logic;
  signal amem5: std_logic;
  signal amem6: std_logic;
  signal amem7: std_logic;
  signal amem8: std_logic;
  signal amem9: std_logic;
  signal amem10: std_logic;
  signal amem11: std_logic;
  signal amem12: std_logic;
  signal amem13: std_logic;
  signal amem14: std_logic;
  signal amem15: std_logic;
  signal amem16: std_logic;
  signal amem17: std_logic;
  signal amem18: std_logic;
  signal amem19: std_logic;
  signal amem20: std_logic;
  signal amem21: std_logic;
  signal amem22: std_logic;
  signal amem23: std_logic;
  signal amem24: std_logic;
  signal amem25: std_logic;
  signal amem26: std_logic;
  signal amem27: std_logic;
  signal amem28: std_logic;
  signal amem29: std_logic;
  signal amem30: std_logic;
  signal amem31: std_logic;
  signal \-amemenb\: std_logic;
  signal amemparity: std_logic;
  signal aparity: std_logic;
  signal aparl: std_logic;
  signal aparm: std_logic;
  signal aparok: std_logic;
  signal \-apass\: std_logic;
  signal apass1: std_logic;
  signal apass2: std_logic;
  signal \-apassenb\: std_logic;
  signal apassenb: std_logic;
  signal \-ape\: std_logic;
  signal \-awpa\: std_logic;
  signal \-awpb\: std_logic;
  signal \-awpc\: std_logic;
  signal \-boot\: std_logic;
  signal \boot.trap\: std_logic;
  signal \-boot1\: std_logic;
  signal \-boot2\: std_logic;
  signal \bottom.1k\: std_logic;
  signal \bus.power.reset l\: std_logic;
  signal \-bus.reset\: std_logic;
  signal \-busint.lm.reset\: std_logic;
  signal \-cin0\: std_logic;
  signal \-cin4\: std_logic;
  signal \-cin8\: std_logic;
  signal \-cin12\: std_logic;
  signal \-cin16\: std_logic;
  signal \-cin20\: std_logic;
  signal \-cin24\: std_logic;
  signal \-cin28\: std_logic;
  signal \-cin32\: std_logic;
  signal \-clk0\: std_logic;
  signal \-clk1\: std_logic;
  signal clk1: std_logic;
  signal clk2: std_logic;
  signal clk3: std_logic;
  signal clk4: std_logic;
  signal clk5: std_logic;
  signal \-clk5\: std_logic;
  signal clk1a: std_logic;
  signal \-clk2a\: std_logic;
  signal clk2a: std_logic;
  signal clk2b: std_logic;
  signal \-clk2c\: std_logic;
  signal clk2c: std_logic;
  signal \-clk3a\: std_logic;
  signal clk3a: std_logic;
  signal clk3b: std_logic;
  signal clk3c: std_logic;
  signal clk3d: std_logic;
  signal \-clk3d\: std_logic;
  signal clk3e: std_logic;
  signal clk3f: std_logic;
  signal \-clk3g\: std_logic;
  signal \-clk4a\: std_logic;
  signal clk4a: std_logic;
  signal clk4b: std_logic;
  signal clk4c: std_logic;
  signal \-clk4d\: std_logic;
  signal clk4d: std_logic;
  signal \-clk4e\: std_logic;
  signal clk4e: std_logic;
  signal clk4f: std_logic;
  signal clk5a: std_logic;
  signal \-clock reset a\: std_logic;
  signal \-clock reset b\: std_logic;
  signal conds0: std_logic;
  signal conds1: std_logic;
  signal conds2: std_logic;
  signal cyclecompleted: std_logic;
  signal \-dadr0a\: std_logic;
  signal \-dadr0b\: std_logic;
  signal \-dadr0c\: std_logic;
  signal \-dadr1a\: std_logic;
  signal \-dadr1b\: std_logic;
  signal \-dadr1c\: std_logic;
  signal \-dadr2a\: std_logic;
  signal \-dadr2b\: std_logic;
  signal \-dadr2c\: std_logic;
  signal \-dadr3a\: std_logic;
  signal \-dadr3b\: std_logic;
  signal \-dadr3c\: std_logic;
  signal \-dadr4a\: std_logic;
  signal \-dadr4b\: std_logic;
  signal \-dadr4c\: std_logic;
  signal \-dadr5a\: std_logic;
  signal \-dadr5b\: std_logic;
  signal \-dadr5c\: std_logic;
  signal \-dadr6a\: std_logic;
  signal \-dadr6b\: std_logic;
  signal \-dadr6c\: std_logic;
  signal \-dadr7a\: std_logic;
  signal \-dadr7b\: std_logic;
  signal \-dadr7c\: std_logic;
  signal \-dadr8a\: std_logic;
  signal \-dadr8b\: std_logic;
  signal \-dadr8c\: std_logic;
  signal \-dadr9a\: std_logic;
  signal \-dadr9b\: std_logic;
  signal \-dadr9c\: std_logic;
  signal \-dadr10a\: std_logic;
  signal dadr10a: std_logic;
  signal \-dadr10c\: std_logic;
  signal dadr10c: std_logic;
  signal \-dbread\: std_logic;
  signal \-dbwrite\: std_logic;
  signal dc0: std_logic;
  signal dc1: std_logic;
  signal dc2: std_logic;
  signal dc3: std_logic;
  signal dc4: std_logic;
  signal dc5: std_logic;
  signal dc6: std_logic;
  signal dc7: std_logic;
  signal dc8: std_logic;
  signal dc9: std_logic;
  signal dcdrive: std_logic;
  signal dest: std_logic;
  signal destd: std_logic;
  signal \-destimod0\: std_logic;
  signal \-destimod1\: std_logic;
  signal \-destintctl\: std_logic;
  signal \-destlc\: std_logic;
  signal destm: std_logic;
  signal destmd: std_logic;
  signal \-destmdr\: std_logic;
  signal destmdr: std_logic;
  signal \-destmem\: std_logic;
  signal destmem: std_logic;
  signal \-destpdl(p)\: std_logic;
  signal \-destpdl(x)\: std_logic;
  signal \-destpdlp\: std_logic;
  signal \-destpdltop\: std_logic;
  signal \-destpdlx\: std_logic;
  signal \-destspc\: std_logic;
  signal destspc: std_logic;
  signal \-destspcd\: std_logic;
  signal destspcd: std_logic;
  signal \-destvma\: std_logic;
  signal \-dfall\: std_logic;
  signal dispenb: std_logic;
  signal dispwr: std_logic;
  signal \-div\: std_logic;
  signal divaddcond: std_logic;
  signal \-divposlasttime\: std_logic;
  signal divsubcond: std_logic;
  signal \-dmapbenb\: std_logic;
  signal dmask0: std_logic;
  signal dmask1: std_logic;
  signal dmask2: std_logic;
  signal dmask3: std_logic;
  signal dmask4: std_logic;
  signal dmask5: std_logic;
  signal dmask6: std_logic;
  signal dn: std_logic;
  signal \-dp\: std_logic;
  signal dp: std_logic;
  signal dpar: std_logic;
  signal dpareven: std_logic;
  signal \-dparh\: std_logic;
  signal dparl: std_logic;
  signal dparok: std_logic;
  signal dpc0: std_logic;
  signal dpc1: std_logic;
  signal dpc2: std_logic;
  signal dpc3: std_logic;
  signal dpc4: std_logic;
  signal dpc5: std_logic;
  signal dpc6: std_logic;
  signal dpc7: std_logic;
  signal dpc8: std_logic;
  signal dpc9: std_logic;
  signal dpc10: std_logic;
  signal dpc11: std_logic;
  signal dpc12: std_logic;
  signal dpc13: std_logic;
  signal \-dpe\: std_logic;
  signal dpe: std_logic;
  signal \-dr\: std_logic;
  signal dr: std_logic;
  signal \-dwea\: std_logic;
  signal \-dweb\: std_logic;
  signal \-dwec\: std_logic;
  signal eadr0: std_logic;
  signal eadr1: std_logic;
  signal eadr2: std_logic;
  signal eadr3: std_logic;
  signal err: std_logic;
  signal \-errhalt\: std_logic;
  signal errstop: std_logic;
  signal \-funct0\: std_logic;
  signal \-funct1\: std_logic;
  signal \-funct2\: std_logic;
  signal \-funct3\: std_logic;
  signal \-halt\: std_logic;
  signal \-halted\: std_logic;
  signal \-hang\: std_logic;
  signal \have wrong word\: std_logic;
  signal hi1: std_logic;
  signal hi2: std_logic;
  signal hi3: std_logic;
  signal hi4: std_logic;
  signal hi5: std_logic;
  signal hi6: std_logic;
  signal hi7: std_logic;
  signal hi8: std_logic;
  signal hi9: std_logic;
  signal hi10: std_logic;
  signal hi11: std_logic;
  signal hi12: std_logic;
  signal \-higherr\: std_logic;
  signal highok: std_logic;
  signal i0: std_logic;
  signal i1: std_logic;
  signal i2: std_logic;
  signal i3: std_logic;
  signal i4: std_logic;
  signal i5: std_logic;
  signal i6: std_logic;
  signal i7: std_logic;
  signal i8: std_logic;
  signal i9: std_logic;
  signal i10: std_logic;
  signal i11: std_logic;
  signal i12: std_logic;
  signal i13: std_logic;
  signal i14: std_logic;
  signal i15: std_logic;
  signal i16: std_logic;
  signal i17: std_logic;
  signal i18: std_logic;
  signal i19: std_logic;
  signal i20: std_logic;
  signal i21: std_logic;
  signal i22: std_logic;
  signal i23: std_logic;
  signal i24: std_logic;
  signal i25: std_logic;
  signal i26: std_logic;
  signal i27: std_logic;
  signal i28: std_logic;
  signal i29: std_logic;
  signal i30: std_logic;
  signal i31: std_logic;
  signal i32: std_logic;
  signal i33: std_logic;
  signal i34: std_logic;
  signal i35: std_logic;
  signal i36: std_logic;
  signal i37: std_logic;
  signal i38: std_logic;
  signal i39: std_logic;
  signal i40: std_logic;
  signal i41: std_logic;
  signal i42: std_logic;
  signal i43: std_logic;
  signal i44: std_logic;
  signal i45: std_logic;
  signal i46: std_logic;
  signal i47: std_logic;
  signal i48: std_logic;
  signal \-ice0a\: std_logic;
  signal \-ice0b\: std_logic;
  signal \-ice0c\: std_logic;
  signal \-ice0d\: std_logic;
  signal \-ice1a\: std_logic;
  signal \-ice1b\: std_logic;
  signal \-ice1c\: std_logic;
  signal \-ice1d\: std_logic;
  signal \-ice2a\: std_logic;
  signal \-ice2b\: std_logic;
  signal \-ice2c\: std_logic;
  signal \-ice2d\: std_logic;
  signal \-ice3a\: std_logic;
  signal \-ice3b\: std_logic;
  signal \-ice3c\: std_logic;
  signal \-ice3d\: std_logic;
  signal \-idebug\: std_logic;
  signal idebug: std_logic;
  signal \-ifetch\: std_logic;
  signal \-ignpar\: std_logic;
  signal \-ignpopj\: std_logic;
  signal \-ilong\: std_logic;
  signal imod: std_logic;
  signal imodd: std_logic;
  signal \-imodd\: std_logic;
  signal \-inop\: std_logic;
  signal inop: std_logic;
  signal \inst in 2nd or 4th quarter\: std_logic;
  signal \inst in left half\: std_logic;
  signal int: std_logic;
  signal \int.enable\: std_logic;
  signal iob0: std_logic;
  signal iob1: std_logic;
  signal iob2: std_logic;
  signal iob3: std_logic;
  signal iob4: std_logic;
  signal iob5: std_logic;
  signal iob6: std_logic;
  signal iob7: std_logic;
  signal iob8: std_logic;
  signal iob9: std_logic;
  signal iob10: std_logic;
  signal iob11: std_logic;
  signal iob12: std_logic;
  signal iob13: std_logic;
  signal iob14: std_logic;
  signal iob15: std_logic;
  signal iob16: std_logic;
  signal iob17: std_logic;
  signal iob18: std_logic;
  signal iob19: std_logic;
  signal iob20: std_logic;
  signal iob21: std_logic;
  signal iob22: std_logic;
  signal iob23: std_logic;
  signal iob24: std_logic;
  signal iob25: std_logic;
  signal iob26: std_logic;
  signal iob27: std_logic;
  signal iob28: std_logic;
  signal iob29: std_logic;
  signal iob30: std_logic;
  signal iob31: std_logic;
  signal iob32: std_logic;
  signal iob33: std_logic;
  signal iob34: std_logic;
  signal iob35: std_logic;
  signal iob36: std_logic;
  signal iob37: std_logic;
  signal iob38: std_logic;
  signal iob39: std_logic;
  signal iob40: std_logic;
  signal iob41: std_logic;
  signal iob42: std_logic;
  signal iob43: std_logic;
  signal iob44: std_logic;
  signal iob45: std_logic;
  signal iob46: std_logic;
  signal iob47: std_logic;
  signal ipar0: std_logic;
  signal ipar1: std_logic;
  signal ipar2: std_logic;
  signal ipar3: std_logic;
  signal iparity: std_logic;
  signal iparok: std_logic;
  signal ipc0: std_logic;
  signal ipc1: std_logic;
  signal ipc2: std_logic;
  signal ipc3: std_logic;
  signal ipc4: std_logic;
  signal ipc5: std_logic;
  signal ipc6: std_logic;
  signal ipc7: std_logic;
  signal ipc8: std_logic;
  signal ipc9: std_logic;
  signal ipc10: std_logic;
  signal ipc11: std_logic;
  signal ipc12: std_logic;
  signal ipc13: std_logic;
  signal \-ipe\: std_logic;
  signal ipe: std_logic;
  signal \-ipopj\: std_logic;
  signal \-ir0\: std_logic;
  signal ir0: std_logic;
  signal \-ir1\: std_logic;
  signal ir1: std_logic;
  signal \-ir2\: std_logic;
  signal ir2: std_logic;
  signal \-ir3\: std_logic;
  signal ir3: std_logic;
  signal \-ir4\: std_logic;
  signal ir4: std_logic;
  signal ir5: std_logic;
  signal ir6: std_logic;
  signal \-ir6\: std_logic;
  signal ir7: std_logic;
  signal \-ir8\: std_logic;
  signal ir8: std_logic;
  signal ir9: std_logic;
  signal ir10: std_logic;
  signal ir11: std_logic;
  signal \-ir12\: std_logic;
  signal ir12: std_logic;
  signal \-ir13\: std_logic;
  signal ir13: std_logic;
  signal ir14: std_logic;
  signal ir15: std_logic;
  signal ir16: std_logic;
  signal ir17: std_logic;
  signal ir18: std_logic;
  signal ir19: std_logic;
  signal ir20: std_logic;
  signal ir21: std_logic;
  signal ir22: std_logic;
  signal \-ir22\: std_logic;
  signal ir23: std_logic;
  signal ir24: std_logic;
  signal ir25: std_logic;
  signal \-ir25\: std_logic;
  signal ir26: std_logic;
  signal ir27: std_logic;
  signal ir28: std_logic;
  signal ir29: std_logic;
  signal ir30: std_logic;
  signal ir31: std_logic;
  signal \-ir31\: std_logic;
  signal ir32: std_logic;
  signal ir33: std_logic;
  signal ir34: std_logic;
  signal ir35: std_logic;
  signal ir36: std_logic;
  signal ir37: std_logic;
  signal ir38: std_logic;
  signal ir39: std_logic;
  signal ir40: std_logic;
  signal ir41: std_logic;
  signal ir42: std_logic;
  signal ir43: std_logic;
  signal ir44: std_logic;
  signal ir45: std_logic;
  signal ir46: std_logic;
  signal ir47: std_logic;
  signal ir48: std_logic;
  signal ir8b: std_logic;
  signal ir9b: std_logic;
  signal ir12b: std_logic;
  signal ir13b: std_logic;
  signal ir14b: std_logic;
  signal ir15b: std_logic;
  signal ir16b: std_logic;
  signal ir17b: std_logic;
  signal ir18b: std_logic;
  signal ir19b: std_logic;
  signal ir20b: std_logic;
  signal ir21b: std_logic;
  signal ir22b: std_logic;
  signal \-iralu\: std_logic;
  signal iralu: std_logic;
  signal \-irbyte\: std_logic;
  signal \-irdisp\: std_logic;
  signal irdisp: std_logic;
  signal \-irjump\: std_logic;
  signal irjump: std_logic;
  signal \-iwea\: std_logic;
  signal \-iweb\: std_logic;
  signal \-iwec\: std_logic;
  signal \-iwed\: std_logic;
  signal \-iwee\: std_logic;
  signal \-iwef\: std_logic;
  signal \-iweg\: std_logic;
  signal \-iweh\: std_logic;
  signal \-iwei\: std_logic;
  signal \-iwej\: std_logic;
  signal \-iwek\: std_logic;
  signal \-iwel\: std_logic;
  signal \-iwem\: std_logic;
  signal \-iwen\: std_logic;
  signal \-iweo\: std_logic;
  signal \-iwep\: std_logic;
  signal iwr0: std_logic;
  signal iwr1: std_logic;
  signal iwr2: std_logic;
  signal iwr3: std_logic;
  signal iwr4: std_logic;
  signal iwr5: std_logic;
  signal iwr6: std_logic;
  signal iwr7: std_logic;
  signal iwr8: std_logic;
  signal iwr9: std_logic;
  signal iwr10: std_logic;
  signal iwr11: std_logic;
  signal iwr12: std_logic;
  signal iwr13: std_logic;
  signal iwr14: std_logic;
  signal iwr15: std_logic;
  signal iwr16: std_logic;
  signal iwr17: std_logic;
  signal iwr18: std_logic;
  signal iwr19: std_logic;
  signal iwr20: std_logic;
  signal iwr21: std_logic;
  signal iwr22: std_logic;
  signal iwr23: std_logic;
  signal iwr24: std_logic;
  signal iwr25: std_logic;
  signal iwr26: std_logic;
  signal iwr27: std_logic;
  signal iwr28: std_logic;
  signal iwr29: std_logic;
  signal iwr30: std_logic;
  signal iwr31: std_logic;
  signal iwr32: std_logic;
  signal iwr33: std_logic;
  signal iwr34: std_logic;
  signal iwr35: std_logic;
  signal iwr36: std_logic;
  signal iwr37: std_logic;
  signal iwr38: std_logic;
  signal iwr39: std_logic;
  signal iwr40: std_logic;
  signal iwr41: std_logic;
  signal iwr42: std_logic;
  signal iwr43: std_logic;
  signal iwr44: std_logic;
  signal iwr45: std_logic;
  signal iwr46: std_logic;
  signal iwr47: std_logic;
  signal iwr48: std_logic;
  signal iwrite: std_logic;
  signal \-iwrited\: std_logic;
  signal iwrited: std_logic;
  signal \-iwriteda\: std_logic;
  signal iwriteda: std_logic;
  signal iwritedb: std_logic;
  signal iwritedc: std_logic;
  signal iwritedd: std_logic;
  signal iwrp1: std_logic;
  signal iwrp2: std_logic;
  signal iwrp3: std_logic;
  signal iwrp4: std_logic;
  signal jcalf: std_logic;
  signal \-jcond\: std_logic;
  signal jcond: std_logic;
  signal jfalse: std_logic;
  signal jret: std_logic;
  signal jretf: std_logic;
  signal l0: std_logic;
  signal l1: std_logic;
  signal l2: std_logic;
  signal l3: std_logic;
  signal l4: std_logic;
  signal l5: std_logic;
  signal l6: std_logic;
  signal l7: std_logic;
  signal l8: std_logic;
  signal l9: std_logic;
  signal l10: std_logic;
  signal l11: std_logic;
  signal l12: std_logic;
  signal l13: std_logic;
  signal l14: std_logic;
  signal l15: std_logic;
  signal l16: std_logic;
  signal l17: std_logic;
  signal l18: std_logic;
  signal l19: std_logic;
  signal l20: std_logic;
  signal l21: std_logic;
  signal l22: std_logic;
  signal l23: std_logic;
  signal l24: std_logic;
  signal l25: std_logic;
  signal l26: std_logic;
  signal l27: std_logic;
  signal l28: std_logic;
  signal l29: std_logic;
  signal l30: std_logic;
  signal l31: std_logic;
  signal \last byte in word\: std_logic;
  signal \lc byte mode\: std_logic;
  signal \-lc modifies mrot\: std_logic;
  signal lc0: std_logic;
  signal lc1: std_logic;
  signal lc2: std_logic;
  signal lc3: std_logic;
  signal lc4: std_logic;
  signal lc5: std_logic;
  signal lc6: std_logic;
  signal lc7: std_logic;
  signal lc8: std_logic;
  signal lc9: std_logic;
  signal lc0b: std_logic;
  signal lc10: std_logic;
  signal lc11: std_logic;
  signal lc12: std_logic;
  signal lc13: std_logic;
  signal lc14: std_logic;
  signal lc15: std_logic;
  signal lc16: std_logic;
  signal lc17: std_logic;
  signal lc18: std_logic;
  signal lc19: std_logic;
  signal lc20: std_logic;
  signal lc21: std_logic;
  signal lc22: std_logic;
  signal lc23: std_logic;
  signal lc24: std_logic;
  signal lc25: std_logic;
  signal lca0: std_logic;
  signal lca1: std_logic;
  signal lca2: std_logic;
  signal lca3: std_logic;
  signal \-lcdrive\: std_logic;
  signal lcdrive: std_logic;
  signal \-lcinc\: std_logic;
  signal lcinc: std_logic;
  signal \-lcry3\: std_logic;
  signal lcry3: std_logic;
  signal \-lcry7\: std_logic;
  signal \-lcry11\: std_logic;
  signal \-lcry15\: std_logic;
  signal \-lcry19\: std_logic;
  signal \-lcry23\: std_logic;
  signal \-ldclk\: std_logic;
  signal \-lddbirh\: std_logic;
  signal \-lddbirl\: std_logic;
  signal \-lddbirm\: std_logic;
  signal \-ldmode\: std_logic;
  signal ldmode: std_logic;
  signal \-ldopc\: std_logic;
  signal \-ldstat\: std_logic;
  signal ldstat: std_logic;
  signal \lm drive enb\: std_logic;
  signal \-loadmd\: std_logic;
  signal loadmd: std_logic;
  signal \-lowerhighok\: std_logic;
  signal lparity: std_logic;
  signal \-lparity\: std_logic;
  signal lparl: std_logic;
  signal \-lparm\: std_logic;
  signal \lpc.hold\: std_logic;
  signal \-lpc.hold\: std_logic;
  signal lpc0: std_logic;
  signal lpc1: std_logic;
  signal lpc2: std_logic;
  signal lpc3: std_logic;
  signal lpc4: std_logic;
  signal lpc5: std_logic;
  signal lpc6: std_logic;
  signal lpc7: std_logic;
  signal lpc8: std_logic;
  signal lpc9: std_logic;
  signal lpc10: std_logic;
  signal lpc11: std_logic;
  signal lpc12: std_logic;
  signal lpc13: std_logic;
  signal \-lvmo22\: std_logic;
  signal \-lvmo23\: std_logic;
  signal m0: std_logic;
  signal m1: std_logic;
  signal m2: std_logic;
  signal m3: std_logic;
  signal m4: std_logic;
  signal m5: std_logic;
  signal m6: std_logic;
  signal m7: std_logic;
  signal m8: std_logic;
  signal m9: std_logic;
  signal m10: std_logic;
  signal m11: std_logic;
  signal m12: std_logic;
  signal m13: std_logic;
  signal m14: std_logic;
  signal m15: std_logic;
  signal m16: std_logic;
  signal m17: std_logic;
  signal m18: std_logic;
  signal m19: std_logic;
  signal m20: std_logic;
  signal m21: std_logic;
  signal m22: std_logic;
  signal m23: std_logic;
  signal m24: std_logic;
  signal m25: std_logic;
  signal m26: std_logic;
  signal m27: std_logic;
  signal m28: std_logic;
  signal m29: std_logic;
  signal m30: std_logic;
  signal m31: std_logic;
  signal m31b: std_logic;
  signal machrun: std_logic;
  signal \-machrun\: std_logic;
  signal \-machruna\: std_logic;
  signal \-madr0a\: std_logic;
  signal \-madr0b\: std_logic;
  signal \-madr1a\: std_logic;
  signal \-madr1b\: std_logic;
  signal \-madr2a\: std_logic;
  signal \-madr2b\: std_logic;
  signal \-madr3a\: std_logic;
  signal \-madr3b\: std_logic;
  signal \-madr4a\: std_logic;
  signal \-madr4b\: std_logic;
  signal \-mapdrive\: std_logic;
  signal mapi8: std_logic;
  signal mapi9: std_logic;
  signal mapi10: std_logic;
  signal mapi11: std_logic;
  signal mapi12: std_logic;
  signal mapi13: std_logic;
  signal mapi14: std_logic;
  signal mapi15: std_logic;
  signal mapi16: std_logic;
  signal mapi17: std_logic;
  signal mapi18: std_logic;
  signal mapi19: std_logic;
  signal mapi20: std_logic;
  signal mapi21: std_logic;
  signal mapi22: std_logic;
  signal mapi23: std_logic;
  signal \-mapi23\: std_logic;
  signal \-mapi8a\: std_logic;
  signal \-mapi8b\: std_logic;
  signal \-mapi9a\: std_logic;
  signal \-mapi9b\: std_logic;
  signal \-mapi10a\: std_logic;
  signal \-mapi10b\: std_logic;
  signal \-mapi11a\: std_logic;
  signal \-mapi11b\: std_logic;
  signal \-mapi12a\: std_logic;
  signal \-mapi12b\: std_logic;
  signal mapwr0d: std_logic;
  signal mapwr1d: std_logic;
  signal mbusy: std_logic;
  signal \-mbusy.sync\: std_logic;
  signal \mbusy.sync\: std_logic;
  signal \-mclk0\: std_logic;
  signal \-mclk1\: std_logic;
  signal mclk1: std_logic;
  signal mclk5: std_logic;
  signal \-mclk5\: std_logic;
  signal mclk7: std_logic;
  signal mclk1a: std_logic;
  signal mclk5a: std_logic;
  signal \-md0\: std_logic;
  signal \-md1\: std_logic;
  signal \-md2\: std_logic;
  signal \-md3\: std_logic;
  signal \-md4\: std_logic;
  signal \-md5\: std_logic;
  signal \-md6\: std_logic;
  signal \-md7\: std_logic;
  signal \-md8\: std_logic;
  signal \-md9\: std_logic;
  signal \-md10\: std_logic;
  signal \-md11\: std_logic;
  signal \-md12\: std_logic;
  signal \-md13\: std_logic;
  signal \-md14\: std_logic;
  signal \-md15\: std_logic;
  signal \-md16\: std_logic;
  signal \-md17\: std_logic;
  signal \-md18\: std_logic;
  signal \-md19\: std_logic;
  signal \-md20\: std_logic;
  signal \-md21\: std_logic;
  signal \-md22\: std_logic;
  signal \-md23\: std_logic;
  signal \-md24\: std_logic;
  signal \-md25\: std_logic;
  signal \-md26\: std_logic;
  signal \-md27\: std_logic;
  signal \-md28\: std_logic;
  signal \-md29\: std_logic;
  signal \-md30\: std_logic;
  signal \-md31\: std_logic;
  signal mdclk: std_logic;
  signal \-mddrive\: std_logic;
  signal mdgetspar: std_logic;
  signal mdhaspar: std_logic;
  signal mdpar: std_logic;
  signal mdparerr: std_logic;
  signal mdpareven: std_logic;
  signal mdparl: std_logic;
  signal mdparm: std_logic;
  signal mdparodd: std_logic;
  signal \-mds0\: std_logic;
  signal \-mds1\: std_logic;
  signal \-mds2\: std_logic;
  signal \-mds3\: std_logic;
  signal \-mds4\: std_logic;
  signal \-mds5\: std_logic;
  signal \-mds6\: std_logic;
  signal \-mds7\: std_logic;
  signal \-mds8\: std_logic;
  signal \-mds9\: std_logic;
  signal \-mds10\: std_logic;
  signal \-mds11\: std_logic;
  signal \-mds12\: std_logic;
  signal \-mds13\: std_logic;
  signal \-mds14\: std_logic;
  signal \-mds15\: std_logic;
  signal \-mds16\: std_logic;
  signal \-mds17\: std_logic;
  signal \-mds18\: std_logic;
  signal \-mds19\: std_logic;
  signal \-mds20\: std_logic;
  signal \-mds21\: std_logic;
  signal \-mds22\: std_logic;
  signal \-mds23\: std_logic;
  signal \-mds24\: std_logic;
  signal \-mds25\: std_logic;
  signal \-mds26\: std_logic;
  signal \-mds27\: std_logic;
  signal \-mds28\: std_logic;
  signal \-mds29\: std_logic;
  signal \-mds30\: std_logic;
  signal \-mds31\: std_logic;
  signal mdsela: std_logic;
  signal mdselb: std_logic;
  signal mem0: std_logic;
  signal mem1: std_logic;
  signal mem2: std_logic;
  signal mem3: std_logic;
  signal mem4: std_logic;
  signal mem5: std_logic;
  signal mem6: std_logic;
  signal mem7: std_logic;
  signal mem8: std_logic;
  signal mem9: std_logic;
  signal mem10: std_logic;
  signal mem11: std_logic;
  signal mem12: std_logic;
  signal mem13: std_logic;
  signal mem14: std_logic;
  signal mem15: std_logic;
  signal mem16: std_logic;
  signal mem17: std_logic;
  signal mem18: std_logic;
  signal mem19: std_logic;
  signal mem20: std_logic;
  signal mem21: std_logic;
  signal mem22: std_logic;
  signal mem23: std_logic;
  signal mem24: std_logic;
  signal mem25: std_logic;
  signal mem26: std_logic;
  signal mem27: std_logic;
  signal mem28: std_logic;
  signal mem29: std_logic;
  signal mem30: std_logic;
  signal mem31: std_logic;
  signal \-memack\: std_logic;
  signal \-memdrive.a\: std_logic;
  signal \-memdrive.b\: std_logic;
  signal \-memgrant\: std_logic;
  signal \-memop\: std_logic;
  signal \mempar in\: std_logic;
  signal \mempar out\: std_logic;
  signal \-memparok\: std_logic;
  signal memparok: std_logic;
  signal \-mempe\: std_logic;
  signal \-memprepare\: std_logic;
  signal memprepare: std_logic;
  signal \-memrd\: std_logic;
  signal memrq: std_logic;
  signal \-memrq\: std_logic;
  signal \-memstart\: std_logic;
  signal memstart: std_logic;
  signal \-memwr\: std_logic;
  signal mf0: std_logic;
  signal mf1: std_logic;
  signal mf2: std_logic;
  signal mf3: std_logic;
  signal mf4: std_logic;
  signal mf5: std_logic;
  signal mf6: std_logic;
  signal mf7: std_logic;
  signal mf8: std_logic;
  signal mf9: std_logic;
  signal mf10: std_logic;
  signal mf11: std_logic;
  signal mf12: std_logic;
  signal mf13: std_logic;
  signal mf14: std_logic;
  signal mf15: std_logic;
  signal mf16: std_logic;
  signal mf17: std_logic;
  signal mf18: std_logic;
  signal mf19: std_logic;
  signal mf20: std_logic;
  signal mf21: std_logic;
  signal mf22: std_logic;
  signal mf23: std_logic;
  signal mf24: std_logic;
  signal mf25: std_logic;
  signal mf26: std_logic;
  signal mf27: std_logic;
  signal mf28: std_logic;
  signal mf29: std_logic;
  signal mf30: std_logic;
  signal mf31: std_logic;
  signal \-mfdrive\: std_logic;
  signal mfdrive: std_logic;
  signal mfenb: std_logic;
  signal \-mfinish\: std_logic;
  signal \-mfinishd\: std_logic;
  signal mmem0: std_logic;
  signal mmem1: std_logic;
  signal mmem2: std_logic;
  signal mmem3: std_logic;
  signal mmem4: std_logic;
  signal mmem5: std_logic;
  signal mmem6: std_logic;
  signal mmem7: std_logic;
  signal mmem8: std_logic;
  signal mmem9: std_logic;
  signal mmem10: std_logic;
  signal mmem11: std_logic;
  signal mmem12: std_logic;
  signal mmem13: std_logic;
  signal mmem14: std_logic;
  signal mmem15: std_logic;
  signal mmem16: std_logic;
  signal mmem17: std_logic;
  signal mmem18: std_logic;
  signal mmem19: std_logic;
  signal mmem20: std_logic;
  signal mmem21: std_logic;
  signal mmem22: std_logic;
  signal mmem23: std_logic;
  signal mmem24: std_logic;
  signal mmem25: std_logic;
  signal mmem26: std_logic;
  signal mmem27: std_logic;
  signal mmem28: std_logic;
  signal mmem29: std_logic;
  signal mmem30: std_logic;
  signal mmem31: std_logic;
  signal mmemparity: std_logic;
  signal mmemparok: std_logic;
  signal mpareven: std_logic;
  signal mparity: std_logic;
  signal mparl: std_logic;
  signal mparm: std_logic;
  signal mparodd: std_logic;
  signal \-mpass\: std_logic;
  signal mpass: std_logic;
  signal \-mpassl\: std_logic;
  signal mpassl: std_logic;
  signal \-mpassm\: std_logic;
  signal \-mpe\: std_logic;
  signal \-mr\: std_logic;
  signal msk0: std_logic;
  signal msk1: std_logic;
  signal msk2: std_logic;
  signal msk3: std_logic;
  signal msk4: std_logic;
  signal msk5: std_logic;
  signal msk6: std_logic;
  signal msk7: std_logic;
  signal msk8: std_logic;
  signal msk9: std_logic;
  signal msk10: std_logic;
  signal msk11: std_logic;
  signal msk12: std_logic;
  signal msk13: std_logic;
  signal msk14: std_logic;
  signal msk15: std_logic;
  signal msk16: std_logic;
  signal msk17: std_logic;
  signal msk18: std_logic;
  signal msk19: std_logic;
  signal msk20: std_logic;
  signal msk21: std_logic;
  signal msk22: std_logic;
  signal msk23: std_logic;
  signal msk24: std_logic;
  signal msk25: std_logic;
  signal msk26: std_logic;
  signal msk27: std_logic;
  signal msk28: std_logic;
  signal msk29: std_logic;
  signal msk30: std_logic;
  signal msk31: std_logic;
  signal mskl0: std_logic;
  signal mskl1: std_logic;
  signal mskl2: std_logic;
  signal mskl3: std_logic;
  signal mskl4: std_logic;
  signal mskl3cry: std_logic;
  signal mskr0: std_logic;
  signal mskr1: std_logic;
  signal mskr2: std_logic;
  signal mskr3: std_logic;
  signal mskr4: std_logic;
  signal \-mul\: std_logic;
  signal \-mulnop\: std_logic;
  signal \-mwpa\: std_logic;
  signal \-mwpb\: std_logic;
  signal n: std_logic;
  signal needfetch: std_logic;
  signal \-needfetch\: std_logic;
  signal \-newlc\: std_logic;
  signal newlc: std_logic;
  signal \-newlc.in\: std_logic;
  signal \next.instr\: std_logic;
  signal \next.instrd\: std_logic;
  signal \-nop\: std_logic;
  signal nop: std_logic;
  signal \-nop11\: std_logic;
  signal nop11: std_logic;
  signal \-nopa\: std_logic;
  signal nopa: std_logic;
  signal npc0: std_logic;
  signal npc1: std_logic;
  signal npc2: std_logic;
  signal npc3: std_logic;
  signal npc4: std_logic;
  signal npc5: std_logic;
  signal npc6: std_logic;
  signal npc7: std_logic;
  signal npc8: std_logic;
  signal npc9: std_logic;
  signal npc10: std_logic;
  signal npc11: std_logic;
  signal npc12: std_logic;
  signal npc13: std_logic;
  signal ob0: std_logic;
  signal ob1: std_logic;
  signal ob2: std_logic;
  signal ob3: std_logic;
  signal ob4: std_logic;
  signal ob5: std_logic;
  signal ob6: std_logic;
  signal ob7: std_logic;
  signal ob8: std_logic;
  signal ob9: std_logic;
  signal ob10: std_logic;
  signal ob11: std_logic;
  signal ob12: std_logic;
  signal ob13: std_logic;
  signal ob14: std_logic;
  signal ob15: std_logic;
  signal ob16: std_logic;
  signal ob17: std_logic;
  signal ob18: std_logic;
  signal ob19: std_logic;
  signal ob20: std_logic;
  signal ob21: std_logic;
  signal ob22: std_logic;
  signal ob23: std_logic;
  signal ob24: std_logic;
  signal ob25: std_logic;
  signal ob26: std_logic;
  signal ob27: std_logic;
  signal ob28: std_logic;
  signal ob29: std_logic;
  signal ob30: std_logic;
  signal ob31: std_logic;
  signal opc0: std_logic;
  signal opc1: std_logic;
  signal opc2: std_logic;
  signal opc3: std_logic;
  signal opc4: std_logic;
  signal opc5: std_logic;
  signal opc6: std_logic;
  signal opc7: std_logic;
  signal opc8: std_logic;
  signal opc9: std_logic;
  signal opc10: std_logic;
  signal opc11: std_logic;
  signal opc12: std_logic;
  signal opc13: std_logic;
  signal \-opcclk\: std_logic;
  signal opcclk: std_logic;
  signal opcclka: std_logic;
  signal opcclkb: std_logic;
  signal opcclkc: std_logic;
  signal \-opcdrive\: std_logic;
  signal \-opcinh\: std_logic;
  signal opcinh: std_logic;
  signal opcinha: std_logic;
  signal opcinhb: std_logic;
  signal osel0a: std_logic;
  signal osel0b: std_logic;
  signal osel1a: std_logic;
  signal osel1b: std_logic;
  signal \-parerr\: std_logic;
  signal pc0: std_logic;
  signal pc1: std_logic;
  signal pc2: std_logic;
  signal pc3: std_logic;
  signal pc4: std_logic;
  signal pc5: std_logic;
  signal pc6: std_logic;
  signal pc7: std_logic;
  signal pc8: std_logic;
  signal pc9: std_logic;
  signal pc0a: std_logic;
  signal pc0b: std_logic;
  signal pc0c: std_logic;
  signal pc0d: std_logic;
  signal pc0e: std_logic;
  signal pc0f: std_logic;
  signal pc0g: std_logic;
  signal pc0h: std_logic;
  signal pc0i: std_logic;
  signal pc0j: std_logic;
  signal pc0k: std_logic;
  signal pc0l: std_logic;
  signal pc0m: std_logic;
  signal pc0n: std_logic;
  signal pc0o: std_logic;
  signal pc0p: std_logic;
  signal pc10: std_logic;
  signal pc11: std_logic;
  signal pc12: std_logic;
  signal pc13: std_logic;
  signal pc1a: std_logic;
  signal pc1b: std_logic;
  signal pc1c: std_logic;
  signal pc1d: std_logic;
  signal pc1e: std_logic;
  signal pc1f: std_logic;
  signal pc1g: std_logic;
  signal pc1h: std_logic;
  signal pc1i: std_logic;
  signal pc1j: std_logic;
  signal pc1k: std_logic;
  signal pc1l: std_logic;
  signal pc1m: std_logic;
  signal pc1n: std_logic;
  signal pc1o: std_logic;
  signal pc1p: std_logic;
  signal pc2a: std_logic;
  signal pc2b: std_logic;
  signal pc2c: std_logic;
  signal pc2d: std_logic;
  signal pc2e: std_logic;
  signal pc2f: std_logic;
  signal pc2g: std_logic;
  signal pc2h: std_logic;
  signal pc2i: std_logic;
  signal pc2j: std_logic;
  signal pc2k: std_logic;
  signal pc2l: std_logic;
  signal pc2m: std_logic;
  signal pc2n: std_logic;
  signal pc2o: std_logic;
  signal pc2p: std_logic;
  signal pc3a: std_logic;
  signal pc3b: std_logic;
  signal pc3c: std_logic;
  signal pc3d: std_logic;
  signal pc3e: std_logic;
  signal pc3f: std_logic;
  signal pc3g: std_logic;
  signal pc3h: std_logic;
  signal pc3i: std_logic;
  signal pc3j: std_logic;
  signal pc3k: std_logic;
  signal pc3l: std_logic;
  signal pc3m: std_logic;
  signal pc3n: std_logic;
  signal pc3o: std_logic;
  signal pc3p: std_logic;
  signal pc4a: std_logic;
  signal pc4b: std_logic;
  signal pc4c: std_logic;
  signal pc4d: std_logic;
  signal pc4e: std_logic;
  signal pc4f: std_logic;
  signal pc4g: std_logic;
  signal pc4h: std_logic;
  signal pc4i: std_logic;
  signal pc4j: std_logic;
  signal pc4k: std_logic;
  signal pc4l: std_logic;
  signal pc4m: std_logic;
  signal pc4n: std_logic;
  signal pc4o: std_logic;
  signal pc4p: std_logic;
  signal pc5a: std_logic;
  signal pc5b: std_logic;
  signal pc5c: std_logic;
  signal pc5d: std_logic;
  signal pc5e: std_logic;
  signal pc5f: std_logic;
  signal pc5g: std_logic;
  signal pc5h: std_logic;
  signal pc5i: std_logic;
  signal pc5j: std_logic;
  signal pc5k: std_logic;
  signal pc5l: std_logic;
  signal pc5m: std_logic;
  signal pc5n: std_logic;
  signal pc5o: std_logic;
  signal pc5p: std_logic;
  signal pc6a: std_logic;
  signal pc6b: std_logic;
  signal pc6c: std_logic;
  signal pc6d: std_logic;
  signal pc6e: std_logic;
  signal pc6f: std_logic;
  signal pc6g: std_logic;
  signal pc6h: std_logic;
  signal pc6i: std_logic;
  signal pc6j: std_logic;
  signal pc6k: std_logic;
  signal pc6l: std_logic;
  signal pc6m: std_logic;
  signal pc6n: std_logic;
  signal pc6o: std_logic;
  signal pc6p: std_logic;
  signal pc7a: std_logic;
  signal pc7b: std_logic;
  signal pc7c: std_logic;
  signal pc7d: std_logic;
  signal pc7e: std_logic;
  signal pc7f: std_logic;
  signal pc7g: std_logic;
  signal pc7h: std_logic;
  signal pc7i: std_logic;
  signal pc7j: std_logic;
  signal pc7k: std_logic;
  signal pc7l: std_logic;
  signal pc7m: std_logic;
  signal pc7n: std_logic;
  signal pc7o: std_logic;
  signal pc7p: std_logic;
  signal pc8a: std_logic;
  signal pc8b: std_logic;
  signal pc8c: std_logic;
  signal pc8d: std_logic;
  signal pc8e: std_logic;
  signal pc8f: std_logic;
  signal pc8g: std_logic;
  signal pc8h: std_logic;
  signal pc8i: std_logic;
  signal pc8j: std_logic;
  signal pc8k: std_logic;
  signal pc8l: std_logic;
  signal pc8m: std_logic;
  signal pc8n: std_logic;
  signal pc8o: std_logic;
  signal pc8p: std_logic;
  signal pc9a: std_logic;
  signal pc9b: std_logic;
  signal pc9c: std_logic;
  signal pc9d: std_logic;
  signal pc9e: std_logic;
  signal pc9f: std_logic;
  signal pc9g: std_logic;
  signal pc9h: std_logic;
  signal pc9i: std_logic;
  signal pc9j: std_logic;
  signal pc9k: std_logic;
  signal pc9l: std_logic;
  signal pc9m: std_logic;
  signal pc9n: std_logic;
  signal pc9o: std_logic;
  signal pc9p: std_logic;
  signal pc10a: std_logic;
  signal pc10b: std_logic;
  signal pc10c: std_logic;
  signal pc10d: std_logic;
  signal pc10e: std_logic;
  signal pc10f: std_logic;
  signal pc10g: std_logic;
  signal pc10h: std_logic;
  signal pc10i: std_logic;
  signal pc10j: std_logic;
  signal pc10k: std_logic;
  signal pc10l: std_logic;
  signal pc10m: std_logic;
  signal pc10n: std_logic;
  signal pc10o: std_logic;
  signal pc10p: std_logic;
  signal pc11a: std_logic;
  signal pc11b: std_logic;
  signal pc11c: std_logic;
  signal pc11d: std_logic;
  signal pc11e: std_logic;
  signal pc11f: std_logic;
  signal pc11g: std_logic;
  signal pc11h: std_logic;
  signal pc11i: std_logic;
  signal pc11j: std_logic;
  signal pc11k: std_logic;
  signal pc11l: std_logic;
  signal pc11m: std_logic;
  signal pc11n: std_logic;
  signal pc11o: std_logic;
  signal pc11p: std_logic;
  signal pc12b: std_logic;
  signal \-pc12b\: std_logic;
  signal pc13b: std_logic;
  signal \-pc13b\: std_logic;
  signal \-pcb0\: std_logic;
  signal \-pcb1\: std_logic;
  signal \-pcb2\: std_logic;
  signal \-pcb3\: std_logic;
  signal \-pcb4\: std_logic;
  signal \-pcb5\: std_logic;
  signal \-pcb6\: std_logic;
  signal \-pcb7\: std_logic;
  signal \-pcb8\: std_logic;
  signal \-pcb9\: std_logic;
  signal \-pcb10\: std_logic;
  signal \-pcb11\: std_logic;
  signal \-pcc0\: std_logic;
  signal \-pcc1\: std_logic;
  signal \-pcc2\: std_logic;
  signal \-pcc3\: std_logic;
  signal \-pcc4\: std_logic;
  signal \-pcc5\: std_logic;
  signal \-pcc6\: std_logic;
  signal \-pcc7\: std_logic;
  signal \-pcc8\: std_logic;
  signal \-pcc9\: std_logic;
  signal \-pcc10\: std_logic;
  signal \-pcc11\: std_logic;
  signal pccry3: std_logic;
  signal pccry7: std_logic;
  signal pccry11: std_logic;
  signal pcs0: std_logic;
  signal pcs1: std_logic;
  signal pdl0: std_logic;
  signal pdl1: std_logic;
  signal pdl2: std_logic;
  signal pdl3: std_logic;
  signal pdl4: std_logic;
  signal pdl5: std_logic;
  signal pdl6: std_logic;
  signal pdl7: std_logic;
  signal pdl8: std_logic;
  signal pdl9: std_logic;
  signal pdl10: std_logic;
  signal pdl11: std_logic;
  signal pdl12: std_logic;
  signal pdl13: std_logic;
  signal pdl14: std_logic;
  signal pdl15: std_logic;
  signal pdl16: std_logic;
  signal pdl17: std_logic;
  signal pdl18: std_logic;
  signal pdl19: std_logic;
  signal pdl20: std_logic;
  signal pdl21: std_logic;
  signal pdl22: std_logic;
  signal pdl23: std_logic;
  signal pdl24: std_logic;
  signal pdl25: std_logic;
  signal pdl26: std_logic;
  signal pdl27: std_logic;
  signal pdl28: std_logic;
  signal pdl29: std_logic;
  signal pdl30: std_logic;
  signal pdl31: std_logic;
  signal \-pdla0a\: std_logic;
  signal \-pdla0b\: std_logic;
  signal \-pdla1a\: std_logic;
  signal \-pdla1b\: std_logic;
  signal \-pdla2a\: std_logic;
  signal \-pdla2b\: std_logic;
  signal \-pdla3a\: std_logic;
  signal \-pdla3b\: std_logic;
  signal \-pdla4a\: std_logic;
  signal \-pdla4b\: std_logic;
  signal \-pdla5a\: std_logic;
  signal \-pdla5b\: std_logic;
  signal \-pdla6a\: std_logic;
  signal \-pdla6b\: std_logic;
  signal \-pdla7a\: std_logic;
  signal \-pdla7b\: std_logic;
  signal \-pdla8a\: std_logic;
  signal \-pdla8b\: std_logic;
  signal \-pdla9a\: std_logic;
  signal \-pdla9b\: std_logic;
  signal \-pdlcnt\: std_logic;
  signal \-pdlcry3\: std_logic;
  signal \-pdlcry7\: std_logic;
  signal \-pdldrive\: std_logic;
  signal pdlenb: std_logic;
  signal pdlidx0: std_logic;
  signal pdlidx1: std_logic;
  signal pdlidx2: std_logic;
  signal pdlidx3: std_logic;
  signal pdlidx4: std_logic;
  signal pdlidx5: std_logic;
  signal pdlidx6: std_logic;
  signal pdlidx7: std_logic;
  signal pdlidx8: std_logic;
  signal pdlidx9: std_logic;
  signal \-pdlpa\: std_logic;
  signal pdlparity: std_logic;
  signal pdlparok: std_logic;
  signal \-pdlpb\: std_logic;
  signal \-pdlpe\: std_logic;
  signal pdlptr0: std_logic;
  signal pdlptr1: std_logic;
  signal pdlptr2: std_logic;
  signal pdlptr3: std_logic;
  signal pdlptr4: std_logic;
  signal pdlptr5: std_logic;
  signal pdlptr6: std_logic;
  signal pdlptr7: std_logic;
  signal pdlptr8: std_logic;
  signal pdlptr9: std_logic;
  signal pdlwrite: std_logic;
  signal \-pdlwrited\: std_logic;
  signal pdlwrited: std_logic;
  signal \-pfr\: std_logic;
  signal \-pfw\: std_logic;
  signal \pgf.or.int\: std_logic;
  signal \pgf.or.int.or.sb\: std_logic;
  signal pidrive: std_logic;
  signal \-pma8\: std_logic;
  signal \-pma9\: std_logic;
  signal \-pma10\: std_logic;
  signal \-pma11\: std_logic;
  signal \-pma12\: std_logic;
  signal \-pma13\: std_logic;
  signal \-pma14\: std_logic;
  signal \-pma15\: std_logic;
  signal \-pma16\: std_logic;
  signal \-pma17\: std_logic;
  signal \-pma18\: std_logic;
  signal \-pma19\: std_logic;
  signal \-pma20\: std_logic;
  signal \-pma21\: std_logic;
  signal \-popj\: std_logic;
  signal popj: std_logic;
  signal \-power reset\: std_logic;
  signal \power reset a\: std_logic;
  signal \-ppdrive\: std_logic;
  signal \prog.boot\: std_logic;
  signal \prog.bus.reset\: std_logic;
  signal \-prog.reset\: std_logic;
  signal \prog.unibus.reset\: std_logic;
  signal \-promce0\: std_logic;
  signal \-promce1\: std_logic;
  signal promdisable: std_logic;
  signal \-promdisabled\: std_logic;
  signal promdisabled: std_logic;
  signal \-promenable\: std_logic;
  signal promenable: std_logic;
  signal \-prompc0\: std_logic;
  signal \-prompc1\: std_logic;
  signal \-prompc2\: std_logic;
  signal \-prompc3\: std_logic;
  signal \-prompc4\: std_logic;
  signal \-prompc5\: std_logic;
  signal \-prompc6\: std_logic;
  signal \-prompc7\: std_logic;
  signal \-prompc8\: std_logic;
  signal \-prompc9\: std_logic;
  signal \-pwidx\: std_logic;
  signal pwidx: std_logic;
  signal \-pwpa\: std_logic;
  signal \-pwpb\: std_logic;
  signal \-pwpc\: std_logic;
  signal q0: std_logic;
  signal q1: std_logic;
  signal q2: std_logic;
  signal q3: std_logic;
  signal q4: std_logic;
  signal q5: std_logic;
  signal q6: std_logic;
  signal q7: std_logic;
  signal q8: std_logic;
  signal q9: std_logic;
  signal q10: std_logic;
  signal q11: std_logic;
  signal q12: std_logic;
  signal q13: std_logic;
  signal q14: std_logic;
  signal q15: std_logic;
  signal q16: std_logic;
  signal q17: std_logic;
  signal q18: std_logic;
  signal q19: std_logic;
  signal q20: std_logic;
  signal q21: std_logic;
  signal q22: std_logic;
  signal q23: std_logic;
  signal q24: std_logic;
  signal q25: std_logic;
  signal q26: std_logic;
  signal q27: std_logic;
  signal q28: std_logic;
  signal q29: std_logic;
  signal q30: std_logic;
  signal q31: std_logic;
  signal \-qdrive\: std_logic;
  signal qdrive: std_logic;
  signal qs0: std_logic;
  signal qs1: std_logic;
  signal r0: std_logic;
  signal r1: std_logic;
  signal r2: std_logic;
  signal r3: std_logic;
  signal r4: std_logic;
  signal r5: std_logic;
  signal r6: std_logic;
  signal r7: std_logic;
  signal r8: std_logic;
  signal r9: std_logic;
  signal r10: std_logic;
  signal r11: std_logic;
  signal r12: std_logic;
  signal r13: std_logic;
  signal r14: std_logic;
  signal r15: std_logic;
  signal r16: std_logic;
  signal r17: std_logic;
  signal r18: std_logic;
  signal r19: std_logic;
  signal r20: std_logic;
  signal r21: std_logic;
  signal r22: std_logic;
  signal r23: std_logic;
  signal r24: std_logic;
  signal r25: std_logic;
  signal r26: std_logic;
  signal r27: std_logic;
  signal r28: std_logic;
  signal r29: std_logic;
  signal r30: std_logic;
  signal r31: std_logic;
  signal ramdisable: std_logic;
  signal \rd.in.progress\: std_logic;
  signal rdcyc: std_logic;
  signal \-rdfinish\: std_logic;
  signal \-reset\: std_logic;
  signal reset: std_logic;
  signal reta0: std_logic;
  signal reta1: std_logic;
  signal reta2: std_logic;
  signal reta3: std_logic;
  signal reta4: std_logic;
  signal reta5: std_logic;
  signal reta6: std_logic;
  signal reta7: std_logic;
  signal reta8: std_logic;
  signal reta9: std_logic;
  signal reta10: std_logic;
  signal reta11: std_logic;
  signal reta12: std_logic;
  signal reta13: std_logic;
  signal \-run\: std_logic;
  signal run: std_logic;
  signal s0: std_logic;
  signal s1: std_logic;
  signal \-s4\: std_logic;
  signal s4: std_logic;
  signal s2a: std_logic;
  signal s2b: std_logic;
  signal s3a: std_logic;
  signal s3b: std_logic;
  signal sa0: std_logic;
  signal sa1: std_logic;
  signal sa2: std_logic;
  signal sa3: std_logic;
  signal sa4: std_logic;
  signal sa5: std_logic;
  signal sa6: std_logic;
  signal sa7: std_logic;
  signal sa8: std_logic;
  signal sa9: std_logic;
  signal sa10: std_logic;
  signal sa11: std_logic;
  signal sa12: std_logic;
  signal sa13: std_logic;
  signal sa14: std_logic;
  signal sa15: std_logic;
  signal sa16: std_logic;
  signal sa17: std_logic;
  signal sa18: std_logic;
  signal sa19: std_logic;
  signal sa20: std_logic;
  signal sa21: std_logic;
  signal sa22: std_logic;
  signal sa23: std_logic;
  signal sa24: std_logic;
  signal sa25: std_logic;
  signal sa26: std_logic;
  signal sa27: std_logic;
  signal sa28: std_logic;
  signal sa29: std_logic;
  signal sa30: std_logic;
  signal sa31: std_logic;
  signal \sequence.break\: std_logic;
  signal \set.rd.in.progress\: std_logic;
  signal \-sh3\: std_logic;
  signal \-sh4\: std_logic;
  signal sint: std_logic;
  signal sintr: std_logic;
  signal spc0: std_logic;
  signal spc1: std_logic;
  signal spc2: std_logic;
  signal spc3: std_logic;
  signal spc4: std_logic;
  signal spc5: std_logic;
  signal spc6: std_logic;
  signal spc7: std_logic;
  signal spc8: std_logic;
  signal spc9: std_logic;
  signal spc10: std_logic;
  signal spc11: std_logic;
  signal spc12: std_logic;
  signal spc13: std_logic;
  signal spc14: std_logic;
  signal spc15: std_logic;
  signal spc16: std_logic;
  signal spc17: std_logic;
  signal spc18: std_logic;
  signal spc1a: std_logic;
  signal \-spccry\: std_logic;
  signal \-spcdrive\: std_logic;
  signal spcdrive: std_logic;
  signal spcenb: std_logic;
  signal spcmung: std_logic;
  signal \-spcnt\: std_logic;
  signal spco0: std_logic;
  signal spco1: std_logic;
  signal spco2: std_logic;
  signal spco3: std_logic;
  signal spco4: std_logic;
  signal spco5: std_logic;
  signal spco6: std_logic;
  signal spco7: std_logic;
  signal spco8: std_logic;
  signal spco9: std_logic;
  signal spco10: std_logic;
  signal spco11: std_logic;
  signal spco12: std_logic;
  signal spco13: std_logic;
  signal spco14: std_logic;
  signal spco15: std_logic;
  signal spco16: std_logic;
  signal spco17: std_logic;
  signal spco18: std_logic;
  signal spcopar: std_logic;
  signal spcpar: std_logic;
  signal spcparh: std_logic;
  signal spcparok: std_logic;
  signal \-spcpass\: std_logic;
  signal spcptr0: std_logic;
  signal spcptr1: std_logic;
  signal spcptr2: std_logic;
  signal spcptr3: std_logic;
  signal spcptr4: std_logic;
  signal spcw0: std_logic;
  signal spcw1: std_logic;
  signal spcw2: std_logic;
  signal spcw3: std_logic;
  signal spcw4: std_logic;
  signal spcw5: std_logic;
  signal spcw6: std_logic;
  signal spcw7: std_logic;
  signal spcw8: std_logic;
  signal spcw9: std_logic;
  signal spcw10: std_logic;
  signal spcw11: std_logic;
  signal spcw12: std_logic;
  signal spcw13: std_logic;
  signal spcw14: std_logic;
  signal spcw15: std_logic;
  signal spcw16: std_logic;
  signal spcw17: std_logic;
  signal spcw18: std_logic;
  signal spcwpar: std_logic;
  signal spcwparh: std_logic;
  signal \-spcwparl\: std_logic;
  signal \-spcwpass\: std_logic;
  signal spcwpass: std_logic;
  signal \-spe\: std_logic;
  signal \-specalu\: std_logic;
  signal speed0: std_logic;
  signal speed1: std_logic;
  signal speed0a: std_logic;
  signal speed1a: std_logic;
  signal speedclk: std_logic;
  signal \-spop\: std_logic;
  signal \-spush\: std_logic;
  signal spush: std_logic;
  signal \-spushd\: std_logic;
  signal spushd: std_logic;
  signal \-spy.ah\: std_logic;
  signal \-spy.al\: std_logic;
  signal \-spy.flag1\: std_logic;
  signal \-spy.flag2\: std_logic;
  signal \-spy.irh\: std_logic;
  signal \-spy.irl\: std_logic;
  signal \-spy.irm\: std_logic;
  signal \-spy.mh\: std_logic;
  signal \-spy.ml\: std_logic;
  signal \-spy.obh\: std_logic;
  signal \-spy.obl\: std_logic;
  signal \-spy.opc\: std_logic;
  signal \-spy.pc\: std_logic;
  signal \-spy.sth\: std_logic;
  signal \-spy.stl\: std_logic;
  signal spy0: std_logic;
  signal spy1: std_logic;
  signal spy2: std_logic;
  signal spy3: std_logic;
  signal spy4: std_logic;
  signal spy5: std_logic;
  signal spy6: std_logic;
  signal spy7: std_logic;
  signal spy8: std_logic;
  signal spy9: std_logic;
  signal spy10: std_logic;
  signal spy11: std_logic;
  signal spy12: std_logic;
  signal spy13: std_logic;
  signal spy14: std_logic;
  signal spy15: std_logic;
  signal \-sr\: std_logic;
  signal \-srcdc\: std_logic;
  signal \-srclc\: std_logic;
  signal srclc: std_logic;
  signal srcm: std_logic;
  signal \-srcm\: std_logic;
  signal \-srcmap\: std_logic;
  signal srcmap: std_logic;
  signal \-srcmd\: std_logic;
  signal srcmd: std_logic;
  signal \-srcopc\: std_logic;
  signal \-srcpdlidx\: std_logic;
  signal srcpdlidx: std_logic;
  signal \-srcpdlpop\: std_logic;
  signal \-srcpdlptr\: std_logic;
  signal srcpdlptr: std_logic;
  signal \-srcpdltop\: std_logic;
  signal \-srcq\: std_logic;
  signal srcq: std_logic;
  signal \-srcspc\: std_logic;
  signal \-srcspcpop\: std_logic;
  signal \-srcspcpopreal\: std_logic;
  signal \-srcvma\: std_logic;
  signal srcvma: std_logic;
  signal srun: std_logic;
  signal \-ssdone\: std_logic;
  signal ssdone: std_logic;
  signal sspeed0: std_logic;
  signal sspeed1: std_logic;
  signal sstep: std_logic;
  signal st0: std_logic;
  signal st1: std_logic;
  signal st2: std_logic;
  signal st3: std_logic;
  signal st4: std_logic;
  signal st5: std_logic;
  signal st6: std_logic;
  signal st7: std_logic;
  signal st8: std_logic;
  signal st9: std_logic;
  signal st10: std_logic;
  signal st11: std_logic;
  signal st12: std_logic;
  signal st13: std_logic;
  signal st14: std_logic;
  signal st15: std_logic;
  signal st16: std_logic;
  signal st17: std_logic;
  signal st18: std_logic;
  signal st19: std_logic;
  signal st20: std_logic;
  signal st21: std_logic;
  signal st22: std_logic;
  signal st23: std_logic;
  signal st24: std_logic;
  signal st25: std_logic;
  signal st26: std_logic;
  signal st27: std_logic;
  signal st28: std_logic;
  signal st29: std_logic;
  signal st30: std_logic;
  signal st31: std_logic;
  signal \stat.ovf\: std_logic;
  signal \-statbit\: std_logic;
  signal \-stathalt\: std_logic;
  signal stathenb: std_logic;
  signal statstop: std_logic;
  signal \-stc4\: std_logic;
  signal \-stc8\: std_logic;
  signal \-stc12\: std_logic;
  signal \-stc16\: std_logic;
  signal \-stc20\: std_logic;
  signal \-stc24\: std_logic;
  signal \-stc28\: std_logic;
  signal \-stc32\: std_logic;
  signal \-step\: std_logic;
  signal step: std_logic;
  signal \-swpa\: std_logic;
  signal \-swpb\: std_logic;
  signal tilt0: std_logic;
  signal tilt1: std_logic;
  signal \-tpclk\: std_logic;
  signal tpclk: std_logic;
  signal \-tpr0\: std_logic;
  signal \-tpr5\: std_logic;
  signal \-tpr10\: std_logic;
  signal \-tpr15\: std_logic;
  signal \-tpr20\: std_logic;
  signal \-tpr25\: std_logic;
  signal \-tpr40\: std_logic;
  signal \-tpr60\: std_logic;
  signal \-tpr65\: std_logic;
  signal \-tpr70\: std_logic;
  signal \-tpr75\: std_logic;
  signal \-tpr80\: std_logic;
  signal \-tpr85\: std_logic;
  signal \-tpr100\: std_logic;
  signal \-tpr105\: std_logic;
  signal \-tpr110\: std_logic;
  signal \-tpr115\: std_logic;
  signal \-tpr120\: std_logic;
  signal \-tpr125\: std_logic;
  signal \-tpr140\: std_logic;
  signal \-tpr160\: std_logic;
  signal \-tpr180\: std_logic;
  signal \-tpr200\: std_logic;
  signal \-tpr20a\: std_logic;
  signal \-tpr80a\: std_logic;
  signal \-tpr120a\: std_logic;
  signal \-tprend\: std_logic;
  signal tprend: std_logic;
  signal \-tptse\: std_logic;
  signal tptse: std_logic;
  signal \-tpw10\: std_logic;
  signal \-tpw20\: std_logic;
  signal \-tpw25\: std_logic;
  signal \-tpw30\: std_logic;
  signal \-tpw35\: std_logic;
  signal \-tpw40\: std_logic;
  signal \-tpw45\: std_logic;
  signal \-tpw50\: std_logic;
  signal \-tpw55\: std_logic;
  signal \-tpw60\: std_logic;
  signal \-tpw65\: std_logic;
  signal \-tpw70\: std_logic;
  signal \-tpw75\: std_logic;
  signal \-tpw30a\: std_logic;
  signal \-tpw40a\: std_logic;
  signal tpwp: std_logic;
  signal tpwpiram: std_logic;
  signal \-trap\: std_logic;
  signal trapa: std_logic;
  signal trapb: std_logic;
  signal \-trapenb\: std_logic;
  signal trapenb: std_logic;
  signal \-tse1\: std_logic;
  signal \-tse2\: std_logic;
  signal tse2: std_logic;
  signal \-tse3\: std_logic;
  signal \-tse4\: std_logic;
  signal tse1a: std_logic;
  signal tse1b: std_logic;
  signal tse3a: std_logic;
  signal tse4a: std_logic;
  signal tse4b: std_logic;
  signal \-upperhighok\: std_logic;
  signal \-use.map\: std_logic;
  signal \use.md\: std_logic;
  signal \-v0pe\: std_logic;
  signal \-v1pe\: std_logic;
  signal v0parok: std_logic;
  signal vm0pari: std_logic;
  signal \-vm0wpa\: std_logic;
  signal \-vm0wpb\: std_logic;
  signal \-vm1lpar\: std_logic;
  signal vm1mpar: std_logic;
  signal vm1pari: std_logic;
  signal \-vm1wpa\: std_logic;
  signal \-vm1wpb\: std_logic;
  signal \-vma0\: std_logic;
  signal \-vma1\: std_logic;
  signal \-vma2\: std_logic;
  signal \-vma3\: std_logic;
  signal \-vma4\: std_logic;
  signal \-vma5\: std_logic;
  signal \-vma6\: std_logic;
  signal \-vma7\: std_logic;
  signal \-vma8\: std_logic;
  signal \-vma9\: std_logic;
  signal \-vma10\: std_logic;
  signal \-vma11\: std_logic;
  signal \-vma12\: std_logic;
  signal \-vma13\: std_logic;
  signal \-vma14\: std_logic;
  signal \-vma15\: std_logic;
  signal \-vma16\: std_logic;
  signal \-vma17\: std_logic;
  signal \-vma18\: std_logic;
  signal \-vma19\: std_logic;
  signal \-vma20\: std_logic;
  signal \-vma21\: std_logic;
  signal \-vma22\: std_logic;
  signal \-vma23\: std_logic;
  signal \-vma24\: std_logic;
  signal \-vma25\: std_logic;
  signal \-vma26\: std_logic;
  signal \-vma27\: std_logic;
  signal \-vma28\: std_logic;
  signal \-vma29\: std_logic;
  signal \-vma30\: std_logic;
  signal \-vma31\: std_logic;
  signal \-vmadrive\: std_logic;
  signal \-vmaenb\: std_logic;
  signal \-vmaok\: std_logic;
  signal \-vmap0\: std_logic;
  signal \-vmap1\: std_logic;
  signal \-vmap2\: std_logic;
  signal \-vmap3\: std_logic;
  signal \-vmap4\: std_logic;
  signal vmap0a: std_logic;
  signal vmap0b: std_logic;
  signal vmap1a: std_logic;
  signal vmap1b: std_logic;
  signal vmap2a: std_logic;
  signal vmap2b: std_logic;
  signal vmap3a: std_logic;
  signal vmap3b: std_logic;
  signal vmap4a: std_logic;
  signal vmap4b: std_logic;
  signal \-vmas0\: std_logic;
  signal \-vmas1\: std_logic;
  signal \-vmas2\: std_logic;
  signal \-vmas3\: std_logic;
  signal \-vmas4\: std_logic;
  signal \-vmas5\: std_logic;
  signal \-vmas6\: std_logic;
  signal \-vmas7\: std_logic;
  signal \-vmas8\: std_logic;
  signal \-vmas9\: std_logic;
  signal \-vmas10\: std_logic;
  signal \-vmas11\: std_logic;
  signal \-vmas12\: std_logic;
  signal \-vmas13\: std_logic;
  signal \-vmas14\: std_logic;
  signal \-vmas15\: std_logic;
  signal \-vmas16\: std_logic;
  signal \-vmas17\: std_logic;
  signal \-vmas18\: std_logic;
  signal \-vmas19\: std_logic;
  signal \-vmas20\: std_logic;
  signal \-vmas21\: std_logic;
  signal \-vmas22\: std_logic;
  signal \-vmas23\: std_logic;
  signal \-vmas24\: std_logic;
  signal \-vmas25\: std_logic;
  signal \-vmas26\: std_logic;
  signal \-vmas27\: std_logic;
  signal \-vmas28\: std_logic;
  signal \-vmas29\: std_logic;
  signal \-vmas30\: std_logic;
  signal \-vmas31\: std_logic;
  signal vmasela: std_logic;
  signal vmaselb: std_logic;
  signal \-vmo0\: std_logic;
  signal \-vmo1\: std_logic;
  signal \-vmo2\: std_logic;
  signal \-vmo3\: std_logic;
  signal \-vmo4\: std_logic;
  signal \-vmo5\: std_logic;
  signal \-vmo6\: std_logic;
  signal \-vmo7\: std_logic;
  signal \-vmo8\: std_logic;
  signal \-vmo9\: std_logic;
  signal \-vmo10\: std_logic;
  signal \-vmo11\: std_logic;
  signal \-vmo12\: std_logic;
  signal \-vmo13\: std_logic;
  signal \-vmo14\: std_logic;
  signal \-vmo15\: std_logic;
  signal \-vmo16\: std_logic;
  signal \-vmo17\: std_logic;
  signal vmo18: std_logic;
  signal \-vmo18\: std_logic;
  signal vmo19: std_logic;
  signal \-vmo19\: std_logic;
  signal \-vmo20\: std_logic;
  signal \-vmo21\: std_logic;
  signal \-vmo22\: std_logic;
  signal \-vmo23\: std_logic;
  signal vmopar: std_logic;
  signal vmoparck: std_logic;
  signal vmoparl: std_logic;
  signal vmoparm: std_logic;
  signal vmoparodd: std_logic;
  signal vmoparok: std_logic;
  signal vpari: std_logic;
  signal wadr0: std_logic;
  signal wadr1: std_logic;
  signal wadr2: std_logic;
  signal wadr3: std_logic;
  signal wadr4: std_logic;
  signal wadr5: std_logic;
  signal wadr6: std_logic;
  signal wadr7: std_logic;
  signal wadr8: std_logic;
  signal wadr9: std_logic;
  signal \-wait\: std_logic;
  signal wmap: std_logic;
  signal \-wmap\: std_logic;
  signal wmapd: std_logic;
  signal \-wmapd\: std_logic;
  signal \-wp1\: std_logic;
  signal \-wp2\: std_logic;
  signal wp2: std_logic;
  signal \-wp3\: std_logic;
  signal \-wp4\: std_logic;
  signal \-wp5\: std_logic;
  signal wp1a: std_logic;
  signal wp1b: std_logic;
  signal wp3a: std_logic;
  signal wp4a: std_logic;
  signal wp4b: std_logic;
  signal wp4c: std_logic;
  signal wp5a: std_logic;
  signal wp5b: std_logic;
  signal wp5c: std_logic;
  signal wp5d: std_logic;
  signal wpc0: std_logic;
  signal wpc1: std_logic;
  signal wpc2: std_logic;
  signal wpc3: std_logic;
  signal wpc4: std_logic;
  signal wpc5: std_logic;
  signal wpc6: std_logic;
  signal wpc7: std_logic;
  signal wpc8: std_logic;
  signal wpc9: std_logic;
  signal wpc10: std_logic;
  signal wpc11: std_logic;
  signal wpc12: std_logic;
  signal wpc13: std_logic;
  signal wrcyc: std_logic;
  signal xout3: std_logic;
  signal xout7: std_logic;
  signal xout11: std_logic;
  signal xout15: std_logic;
  signal xout19: std_logic;
  signal xout23: std_logic;
  signal xout27: std_logic;
  signal xout31: std_logic;
  signal xx0: std_logic;
  signal xx1: std_logic;
  signal yout3: std_logic;
  signal yout7: std_logic;
  signal yout11: std_logic;
  signal yout15: std_logic;
  signal yout19: std_logic;
  signal yout23: std_logic;
  signal yout27: std_logic;
  signal yout31: std_logic;
  signal yy0: std_logic;
  signal yy1: std_logic;
  signal zero16: std_logic;
  signal \zero12.drive\: std_logic;
  signal \-zero16.drive\: std_logic;
  signal \zero16.drive\: std_logic;
begin
  cadr_actl_inst: cadr_actl port map (
      -- in ports
    clk3d => clk3d,
    clk3e => clk3e,
    dest => dest,
    destm => destm,
    hi3 => hi3,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    \-reset\ => \-reset\,
    tse3a => tse3a,
    tse4a => tse4a,
    wp3a => wp3a,
      -- out ports
    \-aadr0a\ => \-aadr0a\,
    \-aadr0b\ => \-aadr0b\,
    \-aadr1a\ => \-aadr1a\,
    \-aadr1b\ => \-aadr1b\,
    \-aadr2a\ => \-aadr2a\,
    \-aadr2b\ => \-aadr2b\,
    \-aadr3a\ => \-aadr3a\,
    \-aadr3b\ => \-aadr3b\,
    \-aadr4a\ => \-aadr4a\,
    \-aadr4b\ => \-aadr4b\,
    \-aadr5a\ => \-aadr5a\,
    \-aadr5b\ => \-aadr5b\,
    \-aadr6a\ => \-aadr6a\,
    \-aadr6b\ => \-aadr6b\,
    \-aadr7a\ => \-aadr7a\,
    \-aadr7b\ => \-aadr7b\,
    \-aadr8a\ => \-aadr8a\,
    \-aadr8b\ => \-aadr8b\,
    \-aadr9a\ => \-aadr9a\,
    \-aadr9b\ => \-aadr9b\,
    \-amemenb\ => \-amemenb\,
    \-apass\ => \-apass\,
    apass1 => apass1,
    apass2 => apass2,
    \-apassenb\ => \-apassenb\,
    apassenb => apassenb,
    \-awpa\ => \-awpa\,
    \-awpb\ => \-awpb\,
    \-awpc\ => \-awpc\,
    destd => destd,
    destmd => destmd,
    wadr0 => wadr0,
    wadr1 => wadr1,
    wadr2 => wadr2,
    wadr3 => wadr3,
    wadr4 => wadr4,
    wadr5 => wadr5,
    wadr6 => wadr6,
    wadr7 => wadr7,
    wadr8 => wadr8,
    wadr9 => wadr9
  );
  cadr_alatch_inst: cadr_alatch port map (
      -- in ports
    amem0 => amem0,
    amem1 => amem1,
    amem2 => amem2,
    amem3 => amem3,
    amem4 => amem4,
    amem5 => amem5,
    amem6 => amem6,
    amem7 => amem7,
    amem8 => amem8,
    amem9 => amem9,
    amem10 => amem10,
    amem11 => amem11,
    amem12 => amem12,
    amem13 => amem13,
    amem14 => amem14,
    amem15 => amem15,
    amem16 => amem16,
    amem17 => amem17,
    amem18 => amem18,
    amem19 => amem19,
    amem20 => amem20,
    amem21 => amem21,
    amem22 => amem22,
    amem23 => amem23,
    amem24 => amem24,
    amem25 => amem25,
    amem26 => amem26,
    amem27 => amem27,
    amem28 => amem28,
    amem29 => amem29,
    amem30 => amem30,
    amem31 => amem31,
    \-amemenb\ => \-amemenb\,
    amemparity => amemparity,
    \-apassenb\ => \-apassenb\,
    apassenb => apassenb,
    clk3e => clk3e,
    hi5 => hi5,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
      -- out ports
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    a31b => a31b,
    aparity => aparity
  );
  cadr_alu0_inst: cadr_alu0 port map (
      -- in ports
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    aluf0b => aluf0b,
    aluf1b => aluf1b,
    aluf2b => aluf2b,
    aluf3b => aluf3b,
    alumode => alumode,
    \-cin0\ => \-cin0\,
    \-cin4\ => \-cin4\,
    \-cin8\ => \-cin8\,
    \-cin12\ => \-cin12\,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
      -- out ports
    \a=m\ => \a=m\,
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    xout3 => xout3,
    xout7 => xout7,
    xout11 => xout11,
    xout15 => xout15,
    yout3 => yout3,
    yout7 => yout7,
    yout11 => yout11,
    yout15 => yout15
  );
  cadr_alu1_inst: cadr_alu1 port map (
      -- in ports
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    a31b => a31b,
    aluf0a => aluf0a,
    aluf1a => aluf1a,
    aluf2a => aluf2a,
    aluf3a => aluf3a,
    alumode => alumode,
    \-cin16\ => \-cin16\,
    \-cin20\ => \-cin20\,
    \-cin24\ => \-cin24\,
    \-cin28\ => \-cin28\,
    \-cin32\ => \-cin32\,
    hi12 => hi12,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
      -- out ports
    \a=m\ => \a=m\,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    alu31 => alu31,
    alu32 => alu32,
    m31b => m31b,
    xout19 => xout19,
    xout23 => xout23,
    xout27 => xout27,
    xout31 => xout31,
    yout19 => yout19,
    yout23 => yout23,
    yout27 => yout27,
    yout31 => yout31
  );
  cadr_aluc4_inst: cadr_aluc4 port map (
      -- in ports
    a31a => a31a,
    a31b => a31b,
    \-div\ => \-div\,
    hi12 => hi12,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    \-ir12\ => \-ir12\,
    \-ir13\ => \-ir13\,
    \-iralu\ => \-iralu\,
    \-irjump\ => \-irjump\,
    irjump => irjump,
    \-mul\ => \-mul\,
    q0 => q0,
    xout3 => xout3,
    xout7 => xout7,
    xout11 => xout11,
    xout19 => xout19,
    xout23 => xout23,
    xout27 => xout27,
    yout3 => yout3,
    yout7 => yout7,
    yout11 => yout11,
    yout19 => yout19,
    yout23 => yout23,
    yout27 => yout27,
      -- out ports
    \-a31\ => \-a31\,
    aluadd => aluadd,
    \-aluf0\ => \-aluf0\,
    \-aluf1\ => \-aluf1\,
    \-aluf2\ => \-aluf2\,
    \-aluf3\ => \-aluf3\,
    aluf0a => aluf0a,
    aluf0b => aluf0b,
    aluf1a => aluf1a,
    aluf1b => aluf1b,
    aluf2a => aluf2a,
    aluf2b => aluf2b,
    aluf3a => aluf3a,
    aluf3b => aluf3b,
    \-alumode\ => \-alumode\,
    alumode => alumode,
    alusub => alusub,
    \-cin0\ => \-cin0\,
    \-cin4\ => \-cin4\,
    \-cin8\ => \-cin8\,
    \-cin12\ => \-cin12\,
    \-cin16\ => \-cin16\,
    \-cin20\ => \-cin20\,
    \-cin24\ => \-cin24\,
    \-cin28\ => \-cin28\,
    \-cin32\ => \-cin32\,
    divaddcond => divaddcond,
    \-divposlasttime\ => \-divposlasttime\,
    divsubcond => divsubcond,
    \-ir0\ => \-ir0\,
    \-ir1\ => \-ir1\,
    \-ir2\ => \-ir2\,
    \-ir3\ => \-ir3\,
    \-ir4\ => \-ir4\,
    \-mulnop\ => \-mulnop\,
    osel0a => osel0a,
    osel0b => osel0b,
    osel1a => osel1a,
    osel1b => osel1b,
    xout15 => xout15,
    xout31 => xout31,
    xx0 => xx0,
    xx1 => xx1,
    yout15 => yout15,
    yout31 => yout31,
    yy0 => yy0,
    yy1 => yy1
  );
  cadr_amem0_inst: cadr_amem0 port map (
      -- in ports
    \-aadr0b\ => \-aadr0b\,
    \-aadr1b\ => \-aadr1b\,
    \-aadr2b\ => \-aadr2b\,
    \-aadr3b\ => \-aadr3b\,
    \-aadr4b\ => \-aadr4b\,
    \-aadr5b\ => \-aadr5b\,
    \-aadr6b\ => \-aadr6b\,
    \-aadr7b\ => \-aadr7b\,
    \-aadr8b\ => \-aadr8b\,
    \-aadr9b\ => \-aadr9b\,
    \-awpa\ => \-awpa\,
    \-awpb\ => \-awpb\,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
      -- out ports
    amem16 => amem16,
    amem17 => amem17,
    amem18 => amem18,
    amem19 => amem19,
    amem20 => amem20,
    amem21 => amem21,
    amem22 => amem22,
    amem23 => amem23,
    amem24 => amem24,
    amem25 => amem25,
    amem26 => amem26,
    amem27 => amem27,
    amem28 => amem28,
    amem29 => amem29,
    amem30 => amem30,
    amem31 => amem31,
    amemparity => amemparity
  );
  cadr_amem1_inst: cadr_amem1 port map (
      -- in ports
    \-aadr0a\ => \-aadr0a\,
    \-aadr1a\ => \-aadr1a\,
    \-aadr2a\ => \-aadr2a\,
    \-aadr3a\ => \-aadr3a\,
    \-aadr4a\ => \-aadr4a\,
    \-aadr5a\ => \-aadr5a\,
    \-aadr6a\ => \-aadr6a\,
    \-aadr7a\ => \-aadr7a\,
    \-aadr8a\ => \-aadr8a\,
    \-aadr9a\ => \-aadr9a\,
    \-awpb\ => \-awpb\,
    \-awpc\ => \-awpc\,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
      -- out ports
    amem0 => amem0,
    amem1 => amem1,
    amem2 => amem2,
    amem3 => amem3,
    amem4 => amem4,
    amem5 => amem5,
    amem6 => amem6,
    amem7 => amem7,
    amem8 => amem8,
    amem9 => amem9,
    amem10 => amem10,
    amem11 => amem11,
    amem12 => amem12,
    amem13 => amem13,
    amem14 => amem14,
    amem15 => amem15
  );
  cadr_apar_inst: cadr_apar port map (
      -- in ports
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31b => a31b,
    aparity => aparity,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    mparity => mparity,
    pdlenb => pdlenb,
    srcm => srcm,
      -- out ports
    aparl => aparl,
    aparm => aparm,
    aparok => aparok,
    mmemparok => mmemparok,
    mpareven => mpareven,
    mparl => mparl,
    mparm => mparm,
    mparodd => mparodd,
    pdlparok => pdlparok
  );
  cadr_bcterm_inst: cadr_bcterm port map (
      -- out ports
    \-ignpar\ => \-ignpar\,
    int => int,
    \-loadmd\ => \-loadmd\,
    mem0 => mem0,
    mem1 => mem1,
    mem2 => mem2,
    mem3 => mem3,
    mem4 => mem4,
    mem5 => mem5,
    mem6 => mem6,
    mem7 => mem7,
    mem8 => mem8,
    mem9 => mem9,
    mem10 => mem10,
    mem11 => mem11,
    mem12 => mem12,
    mem13 => mem13,
    mem14 => mem14,
    mem15 => mem15,
    mem16 => mem16,
    mem17 => mem17,
    mem18 => mem18,
    mem19 => mem19,
    mem20 => mem20,
    mem21 => mem21,
    mem22 => mem22,
    mem23 => mem23,
    mem24 => mem24,
    mem25 => mem25,
    mem26 => mem26,
    mem27 => mem27,
    mem28 => mem28,
    mem29 => mem29,
    mem30 => mem30,
    mem31 => mem31,
    \-memack\ => \-memack\,
    \-memgrant\ => \-memgrant\,
    \mempar in\ => \mempar in\
  );
  cadr_clock1_inst: cadr_clock1 port map (
      -- in ports
    \-clock reset b\ => \-clock reset b\,
    \-hang\ => \-hang\,
    \-ilong\ => \-ilong\,
    sspeed0 => sspeed0,
    sspeed1 => sspeed1,
      -- out ports
    cyclecompleted => cyclecompleted,
    \-tpr0\ => \-tpr0\,
    \-tpr5\ => \-tpr5\,
    \-tpr10\ => \-tpr10\,
    \-tpr15\ => \-tpr15\,
    \-tpr20\ => \-tpr20\,
    \-tpr25\ => \-tpr25\,
    \-tpr40\ => \-tpr40\,
    \-tpr60\ => \-tpr60\,
    \-tpr65\ => \-tpr65\,
    \-tpr70\ => \-tpr70\,
    \-tpr75\ => \-tpr75\,
    \-tpr80\ => \-tpr80\,
    \-tpr85\ => \-tpr85\,
    \-tpr100\ => \-tpr100\,
    \-tpr105\ => \-tpr105\,
    \-tpr110\ => \-tpr110\,
    \-tpr115\ => \-tpr115\,
    \-tpr120\ => \-tpr120\,
    \-tpr125\ => \-tpr125\,
    \-tpr140\ => \-tpr140\,
    \-tpr160\ => \-tpr160\,
    \-tpr180\ => \-tpr180\,
    \-tpr200\ => \-tpr200\,
    \-tpr20a\ => \-tpr20a\,
    \-tpr80a\ => \-tpr80a\,
    \-tpr120a\ => \-tpr120a\,
    \-tprend\ => \-tprend\,
    tprend => tprend,
    \-tpw10\ => \-tpw10\,
    \-tpw20\ => \-tpw20\,
    \-tpw25\ => \-tpw25\,
    \-tpw30\ => \-tpw30\,
    \-tpw35\ => \-tpw35\,
    \-tpw40\ => \-tpw40\,
    \-tpw45\ => \-tpw45\,
    \-tpw50\ => \-tpw50\,
    \-tpw55\ => \-tpw55\,
    \-tpw60\ => \-tpw60\,
    \-tpw65\ => \-tpw65\,
    \-tpw70\ => \-tpw70\,
    \-tpw75\ => \-tpw75\,
    \-tpw30a\ => \-tpw30a\,
    \-tpw40a\ => \-tpw40a\
  );
  cadr_clock2_inst: cadr_clock2 port map (
      -- in ports
    \-clock reset b\ => \-clock reset b\,
    hi1 => hi1,
    machrun => machrun,
    \-machruna\ => \-machruna\,
    \-tpr0\ => \-tpr0\,
    \-tpr5\ => \-tpr5\,
    \-tpr25\ => \-tpr25\,
    \-tprend\ => \-tprend\,
    \-tpw30\ => \-tpw30\,
    \-tpw45\ => \-tpw45\,
    \-tpw70\ => \-tpw70\,
      -- out ports
    \-clk0\ => \-clk0\,
    clk1 => clk1,
    clk2 => clk2,
    clk3 => clk3,
    clk4 => clk4,
    clk5 => clk5,
    \-mclk0\ => \-mclk0\,
    mclk1 => mclk1,
    mclk5 => mclk5,
    mclk7 => mclk7,
    \-tpclk\ => \-tpclk\,
    tpclk => tpclk,
    \-tptse\ => \-tptse\,
    tptse => tptse,
    tpwp => tpwp,
    tpwpiram => tpwpiram,
    \-tse1\ => \-tse1\,
    \-tse2\ => \-tse2\,
    \-tse3\ => \-tse3\,
    \-tse4\ => \-tse4\,
    \-wp1\ => \-wp1\,
    \-wp2\ => \-wp2\,
    \-wp3\ => \-wp3\,
    \-wp4\ => \-wp4\,
    \-wp5\ => \-wp5\
  );
  cadr_clockd_inst: cadr_clockd port map (
      -- in ports
    clk1 => clk1,
    clk2 => clk2,
    clk3 => clk3,
    clk4 => clk4,
    hi1 => hi1,
    hi2 => hi2,
    hi3 => hi3,
    hi4 => hi4,
    hi5 => hi5,
    hi6 => hi6,
    hi7 => hi7,
    hi8 => hi8,
    hi9 => hi9,
    hi10 => hi10,
    hi11 => hi11,
    hi12 => hi12,
    lcry3 => lcry3,
    mclk1 => mclk1,
    reset => reset,
    \-srcpdlidx\ => \-srcpdlidx\,
    \-srcpdlptr\ => \-srcpdlptr\,
    \-tse1\ => \-tse1\,
    \-tse2\ => \-tse2\,
    \-tse3\ => \-tse3\,
    \-tse4\ => \-tse4\,
    \-wp1\ => \-wp1\,
    \-wp2\ => \-wp2\,
    \-wp3\ => \-wp3\,
    \-wp4\ => \-wp4\,
      -- out ports
    \-clk1\ => \-clk1\,
    clk1a => clk1a,
    \-clk2a\ => \-clk2a\,
    clk2a => clk2a,
    clk2b => clk2b,
    \-clk2c\ => \-clk2c\,
    clk2c => clk2c,
    \-clk3a\ => \-clk3a\,
    clk3a => clk3a,
    clk3b => clk3b,
    clk3c => clk3c,
    \-clk3d\ => \-clk3d\,
    clk3d => clk3d,
    clk3e => clk3e,
    clk3f => clk3f,
    \-clk3g\ => \-clk3g\,
    \-clk4a\ => \-clk4a\,
    clk4a => clk4a,
    clk4b => clk4b,
    clk4c => clk4c,
    \-clk4d\ => \-clk4d\,
    clk4d => clk4d,
    \-clk4e\ => \-clk4e\,
    clk4e => clk4e,
    clk4f => clk4f,
    \-lcry3\ => \-lcry3\,
    \-mclk1\ => \-mclk1\,
    mclk1a => mclk1a,
    \-reset\ => \-reset\,
    srcpdlidx => srcpdlidx,
    srcpdlptr => srcpdlptr,
    tse2 => tse2,
    tse1a => tse1a,
    tse1b => tse1b,
    tse3a => tse3a,
    tse4a => tse4a,
    tse4b => tse4b,
    \-upperhighok\ => \-upperhighok\,
    wp2 => wp2,
    wp1a => wp1a,
    wp1b => wp1b,
    wp3a => wp3a,
    wp4a => wp4a,
    wp4b => wp4b,
    wp4c => wp4c
  );
  cadr_contrl_inst: cadr_contrl port map (
      -- in ports
    clk3c => clk3c,
    dp => dp,
    dr => dr,
    \-funct2\ => \-funct2\,
    hi4 => hi4,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir42 => ir42,
    \-irdisp\ => \-irdisp\,
    irdisp => irdisp,
    irjump => irjump,
    \-jcond\ => \-jcond\,
    jcond => jcond,
    \-nop11\ => \-nop11\,
    \-reset\ => \-reset\,
    \-srcspc\ => \-srcspc\,
    \-srcspcpop\ => \-srcspcpop\,
    \-trap\ => \-trap\,
    tse3a => tse3a,
    wp4c => wp4c,
      -- out ports
    \-destspc\ => \-destspc\,
    destspc => destspc,
    \-destspcd\ => \-destspcd\,
    destspcd => destspcd,
    \-dfall\ => \-dfall\,
    dispenb => dispenb,
    dn => dn,
    \-dp\ => \-dp\,
    \-dr\ => \-dr\,
    \-ignpopj\ => \-ignpopj\,
    \-inop\ => \-inop\,
    inop => inop,
    \-ipopj\ => \-ipopj\,
    \-ir6\ => \-ir6\,
    \-ir8\ => \-ir8\,
    iwrite => iwrite,
    \-iwrited\ => \-iwrited\,
    iwrited => iwrited,
    jcalf => jcalf,
    jfalse => jfalse,
    jret => jret,
    jretf => jretf,
    n => n,
    \-nop\ => \-nop\,
    nop => nop,
    \-nopa\ => \-nopa\,
    pcs0 => pcs0,
    pcs1 => pcs1,
    \-popj\ => \-popj\,
    popj => popj,
    \-spcdrive\ => \-spcdrive\,
    spcdrive => spcdrive,
    spcenb => spcenb,
    \-spcnt\ => \-spcnt\,
    \-spcpass\ => \-spcpass\,
    \-spcwpass\ => \-spcwpass\,
    spcwpass => spcwpass,
    \-spop\ => \-spop\,
    \-spush\ => \-spush\,
    spush => spush,
    \-spushd\ => \-spushd\,
    spushd => spushd,
    \-srcspcpopreal\ => \-srcspcpopreal\,
    \-swpa\ => \-swpa\,
    \-swpb\ => \-swpb\
  );
  cadr_debug_inst: cadr_debug port map (
      -- in ports
    \-idebug\ => \-idebug\,
    \-lddbirh\ => \-lddbirh\,
    \-lddbirl\ => \-lddbirl\,
    \-lddbirm\ => \-lddbirm\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47
  );
  cadr_dram0_inst: cadr_dram0 port map (
      -- in ports
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    dispwr => dispwr,
    \-dmapbenb\ => \-dmapbenb\,
    dmask0 => dmask0,
    dmask1 => dmask1,
    dmask2 => dmask2,
    dmask3 => dmask3,
    dmask4 => dmask4,
    dmask5 => dmask5,
    dmask6 => dmask6,
    hi4 => hi4,
    hi6 => hi6,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir8b => ir8b,
    ir9b => ir9b,
    ir20b => ir20b,
    ir21b => ir21b,
    ir22b => ir22b,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    vmo18 => vmo18,
    vmo19 => vmo19,
    wp2 => wp2,
      -- out ports
    \-dadr0a\ => \-dadr0a\,
    \-dadr1a\ => \-dadr1a\,
    \-dadr2a\ => \-dadr2a\,
    \-dadr3a\ => \-dadr3a\,
    \-dadr4a\ => \-dadr4a\,
    \-dadr5a\ => \-dadr5a\,
    \-dadr6a\ => \-dadr6a\,
    \-dadr7a\ => \-dadr7a\,
    \-dadr8a\ => \-dadr8a\,
    \-dadr9a\ => \-dadr9a\,
    \-dadr10a\ => \-dadr10a\,
    dadr10a => dadr10a,
    dpc0 => dpc0,
    dpc1 => dpc1,
    dpc2 => dpc2,
    dpc3 => dpc3,
    dpc4 => dpc4,
    dpc5 => dpc5,
    \-dwea\ => \-dwea\,
    ir12b => ir12b,
    ir13b => ir13b,
    ir14b => ir14b,
    ir15b => ir15b,
    ir16b => ir16b,
    ir17b => ir17b,
    ir18b => ir18b,
    ir19b => ir19b
  );
  cadr_dram1_inst: cadr_dram1 port map (
      -- in ports
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    \-dadr10a\ => \-dadr10a\,
    dadr10a => dadr10a,
    \-dadr10c\ => \-dadr10c\,
    dadr10c => dadr10c,
    dispwr => dispwr,
    \-dmapbenb\ => \-dmapbenb\,
    dmask0 => dmask0,
    dmask1 => dmask1,
    dmask2 => dmask2,
    dmask3 => dmask3,
    dmask4 => dmask4,
    dmask5 => dmask5,
    dmask6 => dmask6,
    hi6 => hi6,
    ir8 => ir8,
    ir9 => ir9,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir12b => ir12b,
    ir13b => ir13b,
    ir14b => ir14b,
    ir15b => ir15b,
    ir16b => ir16b,
    ir17b => ir17b,
    ir18b => ir18b,
    ir19b => ir19b,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    wp2 => wp2,
      -- out ports
    \-dadr0b\ => \-dadr0b\,
    \-dadr1b\ => \-dadr1b\,
    \-dadr2b\ => \-dadr2b\,
    \-dadr3b\ => \-dadr3b\,
    \-dadr4b\ => \-dadr4b\,
    \-dadr5b\ => \-dadr5b\,
    \-dadr6b\ => \-dadr6b\,
    \-dadr7b\ => \-dadr7b\,
    \-dadr8b\ => \-dadr8b\,
    \-dadr9b\ => \-dadr9b\,
    dpc6 => dpc6,
    dpc7 => dpc7,
    dpc8 => dpc8,
    dpc9 => dpc9,
    dpc10 => dpc10,
    dpc11 => dpc11,
    \-dweb\ => \-dweb\,
    ir8b => ir8b,
    ir9b => ir9b,
    ir20b => ir20b,
    ir21b => ir21b,
    ir22b => ir22b,
    \-vmo18\ => \-vmo18\,
    vmo18 => vmo18,
    \-vmo19\ => \-vmo19\,
    vmo19 => vmo19
  );
  cadr_dram2_inst: cadr_dram2 port map (
      -- in ports
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    aa16 => aa16,
    aa17 => aa17,
    dispwr => dispwr,
    \-dmapbenb\ => \-dmapbenb\,
    dmask0 => dmask0,
    dmask1 => dmask1,
    dmask2 => dmask2,
    dmask3 => dmask3,
    dmask4 => dmask4,
    dmask5 => dmask5,
    dmask6 => dmask6,
    hi6 => hi6,
    hi11 => hi11,
    ir8b => ir8b,
    ir9b => ir9b,
    ir12b => ir12b,
    ir13b => ir13b,
    ir14b => ir14b,
    ir15b => ir15b,
    ir16b => ir16b,
    ir17b => ir17b,
    ir18b => ir18b,
    ir19b => ir19b,
    ir20b => ir20b,
    ir21b => ir21b,
    ir22b => ir22b,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    vmo18 => vmo18,
    vmo19 => vmo19,
    wp2 => wp2,
      -- out ports
    \-dadr0c\ => \-dadr0c\,
    \-dadr1c\ => \-dadr1c\,
    \-dadr2c\ => \-dadr2c\,
    \-dadr3c\ => \-dadr3c\,
    \-dadr4c\ => \-dadr4c\,
    \-dadr5c\ => \-dadr5c\,
    \-dadr6c\ => \-dadr6c\,
    \-dadr7c\ => \-dadr7c\,
    \-dadr8c\ => \-dadr8c\,
    \-dadr9c\ => \-dadr9c\,
    \-dadr10c\ => \-dadr10c\,
    dadr10c => dadr10c,
    dn => dn,
    dp => dp,
    dpar => dpar,
    dpc12 => dpc12,
    dpc13 => dpc13,
    dr => dr,
    \-dwec\ => \-dwec\
  );
  cadr_dspctl_inst: cadr_dspctl port map (
      -- in ports
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    clk3e => clk3e,
    dispenb => dispenb,
    dn => dn,
    dp => dp,
    dpar => dpar,
    dpc0 => dpc0,
    dpc1 => dpc1,
    dpc2 => dpc2,
    dpc3 => dpc3,
    dpc4 => dpc4,
    dpc5 => dpc5,
    dpc6 => dpc6,
    dpc7 => dpc7,
    dpc8 => dpc8,
    dpc9 => dpc9,
    dpc10 => dpc10,
    dpc11 => dpc11,
    dpc12 => dpc12,
    dpc13 => dpc13,
    dr => dr,
    \-funct2\ => \-funct2\,
    hi4 => hi4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    \-irdisp\ => \-irdisp\,
      -- out ports
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    aa16 => aa16,
    aa17 => aa17,
    dc0 => dc0,
    dc1 => dc1,
    dc2 => dc2,
    dc3 => dc3,
    dc4 => dc4,
    dc5 => dc5,
    dc6 => dc6,
    dc7 => dc7,
    dc8 => dc8,
    dc9 => dc9,
    dispwr => dispwr,
    \-dmapbenb\ => \-dmapbenb\,
    dmask0 => dmask0,
    dmask1 => dmask1,
    dmask2 => dmask2,
    dmask3 => dmask3,
    dmask4 => dmask4,
    dmask5 => dmask5,
    dmask6 => dmask6,
    dpareven => dpareven,
    \-dparh\ => \-dparh\,
    dparl => dparl,
    dparok => dparok
  );
  cadr_flag_inst: cadr_flag port map (
      -- in ports
    \a=m\ => \a=m\,
    alu32 => alu32,
    clk3c => clk3c,
    \-destintctl\ => \-destintctl\,
    hi4 => hi4,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir5 => ir5,
    ir45 => ir45,
    ir46 => ir46,
    \-nopa\ => \-nopa\,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    r0 => r0,
    \-reset\ => \-reset\,
    sintr => sintr,
    \-vmaok\ => \-vmaok\,
      -- out ports
    \-alu32\ => \-alu32\,
    aluneg => aluneg,
    conds0 => conds0,
    conds1 => conds1,
    conds2 => conds2,
    \-ilong\ => \-ilong\,
    \int.enable\ => \int.enable\,
    \-jcond\ => \-jcond\,
    jcond => jcond,
    \lc byte mode\ => \lc byte mode\,
    \pgf.or.int\ => \pgf.or.int\,
    \pgf.or.int.or.sb\ => \pgf.or.int.or.sb\,
    \prog.unibus.reset\ => \prog.unibus.reset\,
    \sequence.break\ => \sequence.break\,
    sint => sint,
    \-statbit\ => \-statbit\
  );
  cadr_ictl_inst: cadr_ictl port map (
      -- in ports
    hi1 => hi1,
    idebug => idebug,
    \-iwrited\ => \-iwrited\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    promdisabled => promdisabled,
    \-wp5\ => \-wp5\,
      -- out ports
    \-ice0a\ => \-ice0a\,
    \-ice0b\ => \-ice0b\,
    \-ice0c\ => \-ice0c\,
    \-ice0d\ => \-ice0d\,
    \-ice1a\ => \-ice1a\,
    \-ice1b\ => \-ice1b\,
    \-ice1c\ => \-ice1c\,
    \-ice1d\ => \-ice1d\,
    \-ice2a\ => \-ice2a\,
    \-ice2b\ => \-ice2b\,
    \-ice2c\ => \-ice2c\,
    \-ice2d\ => \-ice2d\,
    \-ice3a\ => \-ice3a\,
    \-ice3b\ => \-ice3b\,
    \-ice3c\ => \-ice3c\,
    \-ice3d\ => \-ice3d\,
    \-iwea\ => \-iwea\,
    \-iweb\ => \-iweb\,
    \-iwec\ => \-iwec\,
    \-iwed\ => \-iwed\,
    \-iwee\ => \-iwee\,
    \-iwef\ => \-iwef\,
    \-iweg\ => \-iweg\,
    \-iweh\ => \-iweh\,
    \-iwei\ => \-iwei\,
    \-iwej\ => \-iwej\,
    \-iwek\ => \-iwek\,
    \-iwel\ => \-iwel\,
    \-iwem\ => \-iwem\,
    \-iwen\ => \-iwen\,
    \-iweo\ => \-iweo\,
    \-iwep\ => \-iwep\,
    \-iwriteda\ => \-iwriteda\,
    iwriteda => iwriteda,
    iwritedb => iwritedb,
    iwritedc => iwritedc,
    iwritedd => iwritedd,
    \-pc12b\ => \-pc12b\,
    \-pc13b\ => \-pc13b\,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
    \-promdisabled\ => \-promdisabled\,
    ramdisable => ramdisable,
    wp5a => wp5a,
    wp5b => wp5b,
    wp5c => wp5c,
    wp5d => wp5d
  );
  cadr_ior_inst: cadr_ior port map (
      -- in ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
      -- out ports
    iob0 => iob0,
    iob1 => iob1,
    iob2 => iob2,
    iob3 => iob3,
    iob4 => iob4,
    iob5 => iob5,
    iob6 => iob6,
    iob7 => iob7,
    iob8 => iob8,
    iob9 => iob9,
    iob10 => iob10,
    iob11 => iob11,
    iob12 => iob12,
    iob13 => iob13,
    iob14 => iob14,
    iob15 => iob15,
    iob16 => iob16,
    iob17 => iob17,
    iob18 => iob18,
    iob19 => iob19,
    iob20 => iob20,
    iob21 => iob21,
    iob22 => iob22,
    iob23 => iob23,
    iob24 => iob24,
    iob25 => iob25,
    iob26 => iob26,
    iob27 => iob27,
    iob28 => iob28,
    iob29 => iob29,
    iob30 => iob30,
    iob31 => iob31,
    iob32 => iob32,
    iob33 => iob33,
    iob34 => iob34,
    iob35 => iob35,
    iob36 => iob36,
    iob37 => iob37,
    iob38 => iob38,
    iob39 => iob39,
    iob40 => iob40,
    iob41 => iob41,
    iob42 => iob42,
    iob43 => iob43,
    iob44 => iob44,
    iob45 => iob45,
    iob46 => iob46,
    iob47 => iob47
  );
  cadr_ipar_inst: cadr_ipar port map (
      -- in ports
    imodd => imodd,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir10 => ir10,
    ir11 => ir11,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    ir31 => ir31,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    ir42 => ir42,
    ir43 => ir43,
    ir44 => ir44,
    ir45 => ir45,
    ir46 => ir46,
    ir47 => ir47,
    ir48 => ir48,
      -- out ports
    ipar0 => ipar0,
    ipar1 => ipar1,
    ipar2 => ipar2,
    ipar3 => ipar3,
    iparity => iparity,
    iparok => iparok
  );
  cadr_iram00_inst: cadr_iram00 port map (
      -- in ports
    \-ice0a\ => \-ice0a\,
    \-iwea\ => \-iwea\,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    pc0a => pc0a,
    pc1a => pc1a,
    pc2a => pc2a,
    pc3a => pc3a,
    pc4a => pc4a,
    pc5a => pc5a,
    pc6a => pc6a,
    pc7a => pc7a,
    pc8a => pc8a,
    pc9a => pc9a,
    pc10a => pc10a,
    pc11a => pc11a
  );
  cadr_iram01_inst: cadr_iram01 port map (
      -- in ports
    \-ice1a\ => \-ice1a\,
    \-iweb\ => \-iweb\,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    pc0b => pc0b,
    pc1b => pc1b,
    pc2b => pc2b,
    pc3b => pc3b,
    pc4b => pc4b,
    pc5b => pc5b,
    pc6b => pc6b,
    pc7b => pc7b,
    pc8b => pc8b,
    pc9b => pc9b,
    pc10b => pc10b,
    pc11b => pc11b
  );
  cadr_iram02_inst: cadr_iram02 port map (
      -- in ports
    \-ice2a\ => \-ice2a\,
    \-iwec\ => \-iwec\,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    pc0c => pc0c,
    pc1c => pc1c,
    pc2c => pc2c,
    pc3c => pc3c,
    pc4c => pc4c,
    pc5c => pc5c,
    pc6c => pc6c,
    pc7c => pc7c,
    pc8c => pc8c,
    pc9c => pc9c,
    pc10c => pc10c,
    pc11c => pc11c
  );
  cadr_iram03_inst: cadr_iram03 port map (
      -- in ports
    \-ice3a\ => \-ice3a\,
    \-iwed\ => \-iwed\,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    pc0d => pc0d,
    pc1d => pc1d,
    pc2d => pc2d,
    pc3d => pc3d,
    pc4d => pc4d,
    pc5d => pc5d,
    pc6d => pc6d,
    pc7d => pc7d,
    pc8d => pc8d,
    pc9d => pc9d,
    pc10d => pc10d,
    pc11d => pc11d
  );
  cadr_iram10_inst: cadr_iram10 port map (
      -- in ports
    \-ice0b\ => \-ice0b\,
    \-iwee\ => \-iwee\,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    pc0e => pc0e,
    pc1e => pc1e,
    pc2e => pc2e,
    pc3e => pc3e,
    pc4e => pc4e,
    pc5e => pc5e,
    pc6e => pc6e,
    pc7e => pc7e,
    pc8e => pc8e,
    pc9e => pc9e,
    pc10e => pc10e,
    pc11e => pc11e
  );
  cadr_iram11_inst: cadr_iram11 port map (
      -- in ports
    \-ice1b\ => \-ice1b\,
    \-iwef\ => \-iwef\,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    pc0f => pc0f,
    pc1f => pc1f,
    pc2f => pc2f,
    pc3f => pc3f,
    pc4f => pc4f,
    pc5f => pc5f,
    pc6f => pc6f,
    pc7f => pc7f,
    pc8f => pc8f,
    pc9f => pc9f,
    pc10f => pc10f,
    pc11f => pc11f
  );
  cadr_iram12_inst: cadr_iram12 port map (
      -- in ports
    \-ice2b\ => \-ice2b\,
    \-iweg\ => \-iweg\,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    pc0g => pc0g,
    pc1g => pc1g,
    pc2g => pc2g,
    pc3g => pc3g,
    pc4g => pc4g,
    pc5g => pc5g,
    pc6g => pc6g,
    pc7g => pc7g,
    pc8g => pc8g,
    pc9g => pc9g,
    pc10g => pc10g,
    pc11g => pc11g
  );
  cadr_iram13_inst: cadr_iram13 port map (
      -- in ports
    \-ice3b\ => \-ice3b\,
    \-iweh\ => \-iweh\,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    \-pcb0\ => \-pcb0\,
    \-pcb1\ => \-pcb1\,
    \-pcb2\ => \-pcb2\,
    \-pcb3\ => \-pcb3\,
    \-pcb4\ => \-pcb4\,
    \-pcb5\ => \-pcb5\,
    \-pcb6\ => \-pcb6\,
    \-pcb7\ => \-pcb7\,
    \-pcb8\ => \-pcb8\,
    \-pcb9\ => \-pcb9\,
    \-pcb10\ => \-pcb10\,
    \-pcb11\ => \-pcb11\,
      -- out ports
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    pc0h => pc0h,
    pc1h => pc1h,
    pc2h => pc2h,
    pc3h => pc3h,
    pc4h => pc4h,
    pc5h => pc5h,
    pc6h => pc6h,
    pc7h => pc7h,
    pc8h => pc8h,
    pc9h => pc9h,
    pc10h => pc10h,
    pc11h => pc11h
  );
  cadr_iram20_inst: cadr_iram20 port map (
      -- in ports
    \-ice0c\ => \-ice0c\,
    \-iwei\ => \-iwei\,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    pc0i => pc0i,
    pc1i => pc1i,
    pc2i => pc2i,
    pc3i => pc3i,
    pc4i => pc4i,
    pc5i => pc5i,
    pc6i => pc6i,
    pc7i => pc7i,
    pc8i => pc8i,
    pc9i => pc9i,
    pc10i => pc10i,
    pc11i => pc11i
  );
  cadr_iram21_inst: cadr_iram21 port map (
      -- in ports
    \-ice1c\ => \-ice1c\,
    \-iwej\ => \-iwej\,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    pc0j => pc0j,
    pc1j => pc1j,
    pc2j => pc2j,
    pc3j => pc3j,
    pc4j => pc4j,
    pc5j => pc5j,
    pc6j => pc6j,
    pc7j => pc7j,
    pc8j => pc8j,
    pc9j => pc9j,
    pc10j => pc10j,
    pc11j => pc11j
  );
  cadr_iram22_inst: cadr_iram22 port map (
      -- in ports
    \-ice2c\ => \-ice2c\,
    \-iwek\ => \-iwek\,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    pc0k => pc0k,
    pc1k => pc1k,
    pc2k => pc2k,
    pc3k => pc3k,
    pc4k => pc4k,
    pc5k => pc5k,
    pc6k => pc6k,
    pc7k => pc7k,
    pc8k => pc8k,
    pc9k => pc9k,
    pc10k => pc10k,
    pc11k => pc11k
  );
  cadr_iram23_inst: cadr_iram23 port map (
      -- in ports
    \-ice3c\ => \-ice3c\,
    \-iwel\ => \-iwel\,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    pc0l => pc0l,
    pc1l => pc1l,
    pc2l => pc2l,
    pc3l => pc3l,
    pc4l => pc4l,
    pc5l => pc5l,
    pc6l => pc6l,
    pc7l => pc7l,
    pc8l => pc8l,
    pc9l => pc9l,
    pc10l => pc10l,
    pc11l => pc11l
  );
  cadr_iram30_inst: cadr_iram30 port map (
      -- in ports
    \-ice0d\ => \-ice0d\,
    \-iwem\ => \-iwem\,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    pc0m => pc0m,
    pc1m => pc1m,
    pc2m => pc2m,
    pc3m => pc3m,
    pc4m => pc4m,
    pc5m => pc5m,
    pc6m => pc6m,
    pc7m => pc7m,
    pc8m => pc8m,
    pc9m => pc9m,
    pc10m => pc10m,
    pc11m => pc11m
  );
  cadr_iram31_inst: cadr_iram31 port map (
      -- in ports
    \-ice1d\ => \-ice1d\,
    \-iwen\ => \-iwen\,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    pc0n => pc0n,
    pc1n => pc1n,
    pc2n => pc2n,
    pc3n => pc3n,
    pc4n => pc4n,
    pc5n => pc5n,
    pc6n => pc6n,
    pc7n => pc7n,
    pc8n => pc8n,
    pc9n => pc9n,
    pc10n => pc10n,
    pc11n => pc11n
  );
  cadr_iram32_inst: cadr_iram32 port map (
      -- in ports
    \-ice2d\ => \-ice2d\,
    \-iweo\ => \-iweo\,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    pc0o => pc0o,
    pc1o => pc1o,
    pc2o => pc2o,
    pc3o => pc3o,
    pc4o => pc4o,
    pc5o => pc5o,
    pc6o => pc6o,
    pc7o => pc7o,
    pc8o => pc8o,
    pc9o => pc9o,
    pc10o => pc10o,
    pc11o => pc11o
  );
  cadr_iram33_inst: cadr_iram33 port map (
      -- in ports
    \-ice3d\ => \-ice3d\,
    \-iwep\ => \-iwep\,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48,
    \-pcc0\ => \-pcc0\,
    \-pcc1\ => \-pcc1\,
    \-pcc2\ => \-pcc2\,
    \-pcc3\ => \-pcc3\,
    \-pcc4\ => \-pcc4\,
    \-pcc5\ => \-pcc5\,
    \-pcc6\ => \-pcc6\,
    \-pcc7\ => \-pcc7\,
    \-pcc8\ => \-pcc8\,
    \-pcc9\ => \-pcc9\,
    \-pcc10\ => \-pcc10\,
    \-pcc11\ => \-pcc11\,
      -- out ports
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    pc0p => pc0p,
    pc1p => pc1p,
    pc2p => pc2p,
    pc3p => pc3p,
    pc4p => pc4p,
    pc5p => pc5p,
    pc6p => pc6p,
    pc7p => pc7p,
    pc8p => pc8p,
    pc9p => pc9p,
    pc10p => pc10p,
    pc11p => pc11p
  );
  cadr_ireg_inst: cadr_ireg port map (
      -- in ports
    clk3a => clk3a,
    clk3b => clk3b,
    \-destimod0\ => \-destimod0\,
    \-destimod1\ => \-destimod1\,
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    iob0 => iob0,
    iob1 => iob1,
    iob2 => iob2,
    iob3 => iob3,
    iob4 => iob4,
    iob5 => iob5,
    iob6 => iob6,
    iob7 => iob7,
    iob8 => iob8,
    iob9 => iob9,
    iob10 => iob10,
    iob11 => iob11,
    iob12 => iob12,
    iob13 => iob13,
    iob14 => iob14,
    iob15 => iob15,
    iob16 => iob16,
    iob17 => iob17,
    iob18 => iob18,
    iob19 => iob19,
    iob20 => iob20,
    iob21 => iob21,
    iob22 => iob22,
    iob23 => iob23,
    iob24 => iob24,
    iob25 => iob25,
    iob26 => iob26,
    iob27 => iob27,
    iob28 => iob28,
    iob29 => iob29,
    iob30 => iob30,
    iob31 => iob31,
    iob32 => iob32,
    iob33 => iob33,
    iob34 => iob34,
    iob35 => iob35,
    iob36 => iob36,
    iob37 => iob37,
    iob38 => iob38,
    iob39 => iob39,
    iob40 => iob40,
    iob41 => iob41,
    iob42 => iob42,
    iob43 => iob43,
    iob44 => iob44,
    iob45 => iob45,
    iob46 => iob46,
    iob47 => iob47,
      -- out ports
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir10 => ir10,
    ir11 => ir11,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    ir31 => ir31,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    ir42 => ir42,
    ir43 => ir43,
    ir44 => ir44,
    ir45 => ir45,
    ir46 => ir46,
    ir47 => ir47,
    ir48 => ir48
  );
  cadr_iwr_inst: cadr_iwr port map (
      -- in ports
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    clk2c => clk2c,
    clk4c => clk4c,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
      -- out ports
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47
  );
  cadr_iwrpar_inst: cadr_iwrpar port map (
      -- in ports
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
      -- out ports
    iwr48 => iwr48,
    iwrp1 => iwrp1,
    iwrp2 => iwrp2,
    iwrp3 => iwrp3,
    iwrp4 => iwrp4
  );
  cadr_l_inst: cadr_l port map (
      -- in ports
    clk3f => clk3f,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
      -- out ports
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    \-lparity\ => \-lparity\,
    lparity => lparity,
    lparl => lparl,
    \-lparm\ => \-lparm\
  );
  cadr_lc_inst: cadr_lc port map (
      -- in ports
    clk1a => clk1a,
    clk2a => clk2a,
    clk2c => clk2c,
    \-destlc\ => \-destlc\,
    hi11 => hi11,
    \int.enable\ => \int.enable\,
    \lc byte mode\ => \lc byte mode\,
    lc1 => lc1,
    lc2 => lc2,
    lc3 => lc3,
    lc0b => lc0b,
    \-lcry3\ => \-lcry3\,
    needfetch => needfetch,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    \prog.unibus.reset\ => \prog.unibus.reset\,
    \sequence.break\ => \sequence.break\,
    \-srclc\ => \-srclc\,
    tse1a => tse1a,
      -- out ports
    lc4 => lc4,
    lc5 => lc5,
    lc6 => lc6,
    lc7 => lc7,
    lc8 => lc8,
    lc9 => lc9,
    lc10 => lc10,
    lc11 => lc11,
    lc12 => lc12,
    lc13 => lc13,
    lc14 => lc14,
    lc15 => lc15,
    lc16 => lc16,
    lc17 => lc17,
    lc18 => lc18,
    lc19 => lc19,
    lc20 => lc20,
    lc21 => lc21,
    lc22 => lc22,
    lc23 => lc23,
    lc24 => lc24,
    lc25 => lc25,
    \-lcdrive\ => \-lcdrive\,
    lcdrive => lcdrive,
    \-lcry7\ => \-lcry7\,
    \-lcry11\ => \-lcry11\,
    \-lcry15\ => \-lcry15\,
    \-lcry19\ => \-lcry19\,
    \-lcry23\ => \-lcry23\,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    srclc => srclc
  );
  cadr_lcc_inst: cadr_lcc port map (
      -- in ports
    clk2a => clk2a,
    clk3c => clk3c,
    \-destlc\ => \-destlc\,
    int => int,
    \-ir3\ => \-ir3\,
    \-ir4\ => \-ir4\,
    ir10 => ir10,
    ir11 => ir11,
    ir24 => ir24,
    irdisp => irdisp,
    \lc byte mode\ => \lc byte mode\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    \-reset\ => \-reset\,
    spc1 => spc1,
    spc14 => spc14,
    \-spop\ => \-spop\,
    \-srcspcpopreal\ => \-srcspcpopreal\,
      -- out ports
    \have wrong word\ => \have wrong word\,
    \-ifetch\ => \-ifetch\,
    \inst in 2nd or 4th quarter\ => \inst in 2nd or 4th quarter\,
    \inst in left half\ => \inst in left half\,
    \last byte in word\ => \last byte in word\,
    \-lc modifies mrot\ => \-lc modifies mrot\,
    lc0 => lc0,
    lc1 => lc1,
    lc2 => lc2,
    lc3 => lc3,
    lc0b => lc0b,
    lca0 => lca0,
    lca1 => lca1,
    lca2 => lca2,
    lca3 => lca3,
    \-lcinc\ => \-lcinc\,
    lcinc => lcinc,
    lcry3 => lcry3,
    \-needfetch\ => \-needfetch\,
    needfetch => needfetch,
    \-newlc\ => \-newlc\,
    newlc => newlc,
    \-newlc.in\ => \-newlc.in\,
    \next.instr\ => \next.instr\,
    \next.instrd\ => \next.instrd\,
    \-sh3\ => \-sh3\,
    \-sh4\ => \-sh4\,
    sintr => sintr,
    spc1a => spc1a,
    spcmung => spcmung
  );
  cadr_lpc_inst: cadr_lpc port map (
      -- in ports
    clk4b => clk4b,
    hi5 => hi5,
    ir25 => ir25,
    irdisp => irdisp,
    \lpc.hold\ => \lpc.hold\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
      -- out ports
    lpc0 => lpc0,
    lpc1 => lpc1,
    lpc2 => lpc2,
    lpc3 => lpc3,
    lpc4 => lpc4,
    lpc5 => lpc5,
    lpc6 => lpc6,
    lpc7 => lpc7,
    lpc8 => lpc8,
    lpc9 => lpc9,
    lpc10 => lpc10,
    lpc11 => lpc11,
    lpc12 => lpc12,
    lpc13 => lpc13,
    pc0b => pc0b,
    pc1b => pc1b,
    pc2b => pc2b,
    pc3b => pc3b,
    pc4b => pc4b,
    pc5b => pc5b,
    pc6b => pc6b,
    pc7b => pc7b,
    pc8b => pc8b,
    pc9b => pc9b,
    pc10b => pc10b,
    pc11b => pc11b,
    pc12b => pc12b,
    pc13b => pc13b,
    wpc0 => wpc0,
    wpc1 => wpc1,
    wpc2 => wpc2,
    wpc3 => wpc3,
    wpc4 => wpc4,
    wpc5 => wpc5,
    wpc6 => wpc6,
    wpc7 => wpc7,
    wpc8 => wpc8,
    wpc9 => wpc9,
    wpc10 => wpc10,
    wpc11 => wpc11,
    wpc12 => wpc12,
    wpc13 => wpc13
  );
  cadr_mctl_inst: cadr_mctl port map (
      -- in ports
    clk4e => clk4e,
    destmd => destmd,
    hi2 => hi2,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    \-ir31\ => \-ir31\,
    tse4a => tse4a,
    wadr0 => wadr0,
    wadr1 => wadr1,
    wadr2 => wadr2,
    wadr3 => wadr3,
    wadr4 => wadr4,
    wp4b => wp4b,
      -- out ports
    \-madr0a\ => \-madr0a\,
    \-madr0b\ => \-madr0b\,
    \-madr1a\ => \-madr1a\,
    \-madr1b\ => \-madr1b\,
    \-madr2a\ => \-madr2a\,
    \-madr2b\ => \-madr2b\,
    \-madr3a\ => \-madr3a\,
    \-madr3b\ => \-madr3b\,
    \-madr4a\ => \-madr4a\,
    \-madr4b\ => \-madr4b\,
    mmem0 => mmem0,
    mmem1 => mmem1,
    mmem2 => mmem2,
    mmem3 => mmem3,
    mmem4 => mmem4,
    mmem5 => mmem5,
    mmem6 => mmem6,
    mmem7 => mmem7,
    mmem8 => mmem8,
    mmem9 => mmem9,
    mmem10 => mmem10,
    mmem11 => mmem11,
    mmem12 => mmem12,
    mmem13 => mmem13,
    mmem14 => mmem14,
    mmem15 => mmem15,
    mmem16 => mmem16,
    mmem17 => mmem17,
    mmem18 => mmem18,
    mmem19 => mmem19,
    mmem20 => mmem20,
    mmem21 => mmem21,
    mmem22 => mmem22,
    mmem23 => mmem23,
    mmem24 => mmem24,
    mmem25 => mmem25,
    mmem26 => mmem26,
    mmem27 => mmem27,
    mmem28 => mmem28,
    mmem29 => mmem29,
    mmem30 => mmem30,
    mmem31 => mmem31,
    mmemparity => mmemparity,
    \-mpass\ => \-mpass\,
    mpass => mpass,
    \-mpassl\ => \-mpassl\,
    mpassl => mpassl,
    \-mpassm\ => \-mpassm\,
    \-mwpa\ => \-mwpa\,
    \-mwpb\ => \-mwpb\,
    srcm => srcm
  );
  cadr_md_inst: cadr_md port map (
      -- in ports
    \-clk2c\ => \-clk2c\,
    \-destmdr\ => \-destmdr\,
    \-ignpar\ => \-ignpar\,
    \-loadmd\ => \-loadmd\,
    \-mds0\ => \-mds0\,
    \-mds1\ => \-mds1\,
    \-mds2\ => \-mds2\,
    \-mds3\ => \-mds3\,
    \-mds4\ => \-mds4\,
    \-mds5\ => \-mds5\,
    \-mds6\ => \-mds6\,
    \-mds7\ => \-mds7\,
    \-mds8\ => \-mds8\,
    \-mds9\ => \-mds9\,
    \-mds10\ => \-mds10\,
    \-mds11\ => \-mds11\,
    \-mds12\ => \-mds12\,
    \-mds13\ => \-mds13\,
    \-mds14\ => \-mds14\,
    \-mds15\ => \-mds15\,
    \-mds16\ => \-mds16\,
    \-mds17\ => \-mds17\,
    \-mds18\ => \-mds18\,
    \-mds19\ => \-mds19\,
    \-mds20\ => \-mds20\,
    \-mds21\ => \-mds21\,
    \-mds22\ => \-mds22\,
    \-mds23\ => \-mds23\,
    \-mds24\ => \-mds24\,
    \-mds25\ => \-mds25\,
    \-mds26\ => \-mds26\,
    \-mds27\ => \-mds27\,
    \-mds28\ => \-mds28\,
    \-mds29\ => \-mds29\,
    \-mds30\ => \-mds30\,
    \-mds31\ => \-mds31\,
    \mempar in\ => \mempar in\,
    \-srcmd\ => \-srcmd\,
    tse2 => tse2,
      -- out ports
    destmdr => destmdr,
    loadmd => loadmd,
    \-md0\ => \-md0\,
    \-md1\ => \-md1\,
    \-md2\ => \-md2\,
    \-md3\ => \-md3\,
    \-md4\ => \-md4\,
    \-md5\ => \-md5\,
    \-md6\ => \-md6\,
    \-md7\ => \-md7\,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-md24\ => \-md24\,
    \-md25\ => \-md25\,
    \-md26\ => \-md26\,
    \-md27\ => \-md27\,
    \-md28\ => \-md28\,
    \-md29\ => \-md29\,
    \-md30\ => \-md30\,
    \-md31\ => \-md31\,
    mdclk => mdclk,
    \-mddrive\ => \-mddrive\,
    mdgetspar => mdgetspar,
    mdhaspar => mdhaspar,
    mdpar => mdpar,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    srcmd => srcmd
  );
  cadr_mds_inst: cadr_mds port map (
      -- in ports
    hi11 => hi11,
    \-md0\ => \-md0\,
    \-md1\ => \-md1\,
    \-md2\ => \-md2\,
    \-md3\ => \-md3\,
    \-md4\ => \-md4\,
    \-md5\ => \-md5\,
    \-md6\ => \-md6\,
    \-md7\ => \-md7\,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-md24\ => \-md24\,
    \-md25\ => \-md25\,
    \-md26\ => \-md26\,
    \-md27\ => \-md27\,
    \-md28\ => \-md28\,
    \-md29\ => \-md29\,
    \-md30\ => \-md30\,
    \-md31\ => \-md31\,
    mdparodd => mdparodd,
    mdsela => mdsela,
    mdselb => mdselb,
    \-memdrive.a\ => \-memdrive.a\,
    \-memdrive.b\ => \-memdrive.b\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
      -- out ports
    \-mds0\ => \-mds0\,
    \-mds1\ => \-mds1\,
    \-mds2\ => \-mds2\,
    \-mds3\ => \-mds3\,
    \-mds4\ => \-mds4\,
    \-mds5\ => \-mds5\,
    \-mds6\ => \-mds6\,
    \-mds7\ => \-mds7\,
    \-mds8\ => \-mds8\,
    \-mds9\ => \-mds9\,
    \-mds10\ => \-mds10\,
    \-mds11\ => \-mds11\,
    \-mds12\ => \-mds12\,
    \-mds13\ => \-mds13\,
    \-mds14\ => \-mds14\,
    \-mds15\ => \-mds15\,
    \-mds16\ => \-mds16\,
    \-mds17\ => \-mds17\,
    \-mds18\ => \-mds18\,
    \-mds19\ => \-mds19\,
    \-mds20\ => \-mds20\,
    \-mds21\ => \-mds21\,
    \-mds22\ => \-mds22\,
    \-mds23\ => \-mds23\,
    \-mds24\ => \-mds24\,
    \-mds25\ => \-mds25\,
    \-mds26\ => \-mds26\,
    \-mds27\ => \-mds27\,
    \-mds28\ => \-mds28\,
    \-mds29\ => \-mds29\,
    \-mds30\ => \-mds30\,
    \-mds31\ => \-mds31\,
    mem0 => mem0,
    mem1 => mem1,
    mem2 => mem2,
    mem3 => mem3,
    mem4 => mem4,
    mem5 => mem5,
    mem6 => mem6,
    mem7 => mem7,
    mem8 => mem8,
    mem9 => mem9,
    mem10 => mem10,
    mem11 => mem11,
    mem12 => mem12,
    mem13 => mem13,
    mem14 => mem14,
    mem15 => mem15,
    mem16 => mem16,
    mem17 => mem17,
    mem18 => mem18,
    mem19 => mem19,
    mem20 => mem20,
    mem21 => mem21,
    mem22 => mem22,
    mem23 => mem23,
    mem24 => mem24,
    mem25 => mem25,
    mem26 => mem26,
    mem27 => mem27,
    mem28 => mem28,
    mem29 => mem29,
    mem30 => mem30,
    mem31 => mem31,
    \mempar out\ => \mempar out\
  );
  cadr_mf_inst: cadr_mf port map (
      -- in ports
    \-ir31\ => \-ir31\,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    \-mpass\ => \-mpass\,
    pdlenb => pdlenb,
    spcenb => spcenb,
    tse1a => tse1a,
      -- out ports
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    \-mfdrive\ => \-mfdrive\,
    mfdrive => mfdrive,
    mfenb => mfenb,
    \-srcm\ => \-srcm\
  );
  cadr_mlatch_inst: cadr_mlatch port map (
      -- in ports
    clk4a => clk4a,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    mmem2 => mmem2,
    mmem3 => mmem3,
    mmem5 => mmem5,
    mmem7 => mmem7,
    mmem9 => mmem9,
    mmem11 => mmem11,
    mmem13 => mmem13,
    mmem15 => mmem15,
    mmem17 => mmem17,
    mmem19 => mmem19,
    mmem21 => mmem21,
    mmem23 => mmem23,
    mmem25 => mmem25,
    mmem27 => mmem27,
    mmem29 => mmem29,
    mmem31 => mmem31,
    \-mpassl\ => \-mpassl\,
    mpassl => mpassl,
    \-mpassm\ => \-mpassm\,
      -- out ports
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    mmem0 => mmem0,
    mmem1 => mmem1,
    mmem4 => mmem4,
    mmem6 => mmem6,
    mmem8 => mmem8,
    mmem10 => mmem10,
    mmem12 => mmem12,
    mmem14 => mmem14,
    mmem16 => mmem16,
    mmem18 => mmem18,
    mmem20 => mmem20,
    mmem22 => mmem22,
    mmem24 => mmem24,
    mmem26 => mmem26,
    mmem28 => mmem28,
    mmem30 => mmem30,
    mmemparity => mmemparity,
    mparity => mparity
  );
  cadr_mmem_inst: cadr_mmem port map (
      -- in ports
    hi2 => hi2,
    hi3 => hi3,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
    \-madr0a\ => \-madr0a\,
    \-madr0b\ => \-madr0b\,
    \-madr1a\ => \-madr1a\,
    \-madr1b\ => \-madr1b\,
    \-madr2a\ => \-madr2a\,
    \-madr2b\ => \-madr2b\,
    \-madr3a\ => \-madr3a\,
    \-madr3b\ => \-madr3b\,
    \-madr4a\ => \-madr4a\,
    \-madr4b\ => \-madr4b\,
    \-mwpa\ => \-mwpa\,
    \-mwpb\ => \-mwpb\,
      -- out ports
    mmem0 => mmem0,
    mmem1 => mmem1,
    mmem2 => mmem2,
    mmem3 => mmem3,
    mmem4 => mmem4,
    mmem5 => mmem5,
    mmem6 => mmem6,
    mmem7 => mmem7,
    mmem8 => mmem8,
    mmem9 => mmem9,
    mmem10 => mmem10,
    mmem11 => mmem11,
    mmem12 => mmem12,
    mmem13 => mmem13,
    mmem14 => mmem14,
    mmem15 => mmem15,
    mmem16 => mmem16,
    mmem17 => mmem17,
    mmem18 => mmem18,
    mmem19 => mmem19,
    mmem20 => mmem20,
    mmem21 => mmem21,
    mmem22 => mmem22,
    mmem23 => mmem23,
    mmem24 => mmem24,
    mmem25 => mmem25,
    mmem26 => mmem26,
    mmem27 => mmem27,
    mmem28 => mmem28,
    mmem29 => mmem29,
    mmem30 => mmem30,
    mmem31 => mmem31,
    mmemparity => mmemparity
  );
  cadr_mo0_inst: cadr_mo0 port map (
      -- in ports
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    alu16 => alu16,
    msk0 => msk0,
    msk1 => msk1,
    msk2 => msk2,
    msk3 => msk3,
    msk4 => msk4,
    msk5 => msk5,
    msk6 => msk6,
    msk7 => msk7,
    msk8 => msk8,
    msk9 => msk9,
    msk10 => msk10,
    msk11 => msk11,
    msk12 => msk12,
    msk13 => msk13,
    msk14 => msk14,
    msk15 => msk15,
    osel0b => osel0b,
    osel1b => osel1b,
    q31 => q31,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    r7 => r7,
    r8 => r8,
    r9 => r9,
    r10 => r10,
    r11 => r11,
    r12 => r12,
    r13 => r13,
    r14 => r14,
    r15 => r15,
      -- out ports
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15
  );
  cadr_mo1_inst: cadr_mo1 port map (
      -- in ports
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31b => a31b,
    alu15 => alu15,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    alu31 => alu31,
    alu32 => alu32,
    msk16 => msk16,
    msk17 => msk17,
    msk18 => msk18,
    msk19 => msk19,
    msk20 => msk20,
    msk21 => msk21,
    msk22 => msk22,
    msk23 => msk23,
    msk24 => msk24,
    msk25 => msk25,
    msk26 => msk26,
    msk27 => msk27,
    msk28 => msk28,
    msk29 => msk29,
    msk30 => msk30,
    msk31 => msk31,
    osel0a => osel0a,
    osel1a => osel1a,
    r16 => r16,
    r17 => r17,
    r18 => r18,
    r19 => r19,
    r20 => r20,
    r21 => r21,
    r22 => r22,
    r23 => r23,
    r24 => r24,
    r25 => r25,
    r26 => r26,
    r27 => r27,
    r28 => r28,
    r29 => r29,
    r30 => r30,
    r31 => r31,
      -- out ports
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31
  );
  cadr_mskg4_inst: cadr_mskg4 port map (
      -- in ports
    ir12 => ir12,
    ir13 => ir13,
    ir31 => ir31,
    mskl0 => mskl0,
    mskl1 => mskl1,
    mskl2 => mskl2,
    mskl3 => mskl3,
    mskl4 => mskl4,
    mskr0 => mskr0,
    mskr1 => mskr1,
    mskr2 => mskr2,
    mskr3 => mskr3,
    mskr4 => mskr4,
      -- out ports
    \a=m\ => \a=m\,
    \-ir12\ => \-ir12\,
    \-ir13\ => \-ir13\,
    \-ir31\ => \-ir31\,
    msk0 => msk0,
    msk1 => msk1,
    msk2 => msk2,
    msk3 => msk3,
    msk4 => msk4,
    msk5 => msk5,
    msk6 => msk6,
    msk7 => msk7,
    msk8 => msk8,
    msk9 => msk9,
    msk10 => msk10,
    msk11 => msk11,
    msk12 => msk12,
    msk13 => msk13,
    msk14 => msk14,
    msk15 => msk15,
    msk16 => msk16,
    msk17 => msk17,
    msk18 => msk18,
    msk19 => msk19,
    msk20 => msk20,
    msk21 => msk21,
    msk22 => msk22,
    msk23 => msk23,
    msk24 => msk24,
    msk25 => msk25,
    msk26 => msk26,
    msk27 => msk27,
    msk28 => msk28,
    msk29 => msk29,
    msk30 => msk30,
    msk31 => msk31
  );
  cadr_npc_inst: cadr_npc port map (
      -- in ports
    clk4b => clk4b,
    dpc4 => dpc4,
    hi4 => hi4,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    pcs0 => pcs0,
    pcs1 => pcs1,
    spc1a => spc1a,
    trapa => trapa,
    trapb => trapb,
      -- out ports
    dpc0 => dpc0,
    dpc1 => dpc1,
    dpc2 => dpc2,
    dpc3 => dpc3,
    dpc5 => dpc5,
    dpc6 => dpc6,
    dpc7 => dpc7,
    dpc8 => dpc8,
    dpc9 => dpc9,
    dpc10 => dpc10,
    dpc11 => dpc11,
    dpc12 => dpc12,
    dpc13 => dpc13,
    ipc0 => ipc0,
    ipc1 => ipc1,
    ipc2 => ipc2,
    ipc3 => ipc3,
    ipc4 => ipc4,
    ipc5 => ipc5,
    ipc6 => ipc6,
    ipc7 => ipc7,
    ipc8 => ipc8,
    ipc9 => ipc9,
    ipc10 => ipc10,
    ipc11 => ipc11,
    ipc12 => ipc12,
    ipc13 => ipc13,
    npc0 => npc0,
    npc1 => npc1,
    npc2 => npc2,
    npc3 => npc3,
    npc4 => npc4,
    npc5 => npc5,
    npc6 => npc6,
    npc7 => npc7,
    npc8 => npc8,
    npc9 => npc9,
    npc10 => npc10,
    npc11 => npc11,
    npc12 => npc12,
    npc13 => npc13,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    pccry3 => pccry3,
    pccry7 => pccry7,
    pccry11 => pccry11,
    spc0 => spc0,
    spc2 => spc2,
    spc3 => spc3,
    spc4 => spc4,
    spc5 => spc5,
    spc6 => spc6,
    spc7 => spc7,
    spc8 => spc8,
    spc9 => spc9,
    spc10 => spc10,
    spc11 => spc11,
    spc12 => spc12,
    spc13 => spc13
  );
  cadr_olord1_inst: cadr_olord1 port map (
      -- in ports
    \-boot\ => \-boot\,
    \-clock reset a\ => \-clock reset a\,
    \-errhalt\ => \-errhalt\,
    \-ldclk\ => \-ldclk\,
    \-ldmode\ => \-ldmode\,
    \-ldopc\ => \-ldopc\,
    mclk5a => mclk5a,
    \-reset\ => \-reset\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    statstop => statstop,
    \-stc32\ => \-stc32\,
    \-tpr60\ => \-tpr60\,
    \-wait\ => \-wait\,
      -- out ports
    errstop => errstop,
    \-idebug\ => \-idebug\,
    idebug => idebug,
    \-ldstat\ => \-ldstat\,
    ldstat => ldstat,
    \-lpc.hold\ => \-lpc.hold\,
    \lpc.hold\ => \lpc.hold\,
    \-machrun\ => \-machrun\,
    machrun => machrun,
    \-machruna\ => \-machruna\,
    \-nop11\ => \-nop11\,
    nop11 => nop11,
    \-opcclk\ => \-opcclk\,
    opcclk => opcclk,
    \-opcinh\ => \-opcinh\,
    opcinh => opcinh,
    promdisable => promdisable,
    promdisabled => promdisabled,
    \-run\ => \-run\,
    run => run,
    speed0 => speed0,
    speed1 => speed1,
    speed0a => speed0a,
    speed1a => speed1a,
    speedclk => speedclk,
    srun => srun,
    \-ssdone\ => \-ssdone\,
    ssdone => ssdone,
    sspeed0 => sspeed0,
    sspeed1 => sspeed1,
    sstep => sstep,
    \stat.ovf\ => \stat.ovf\,
    \-stathalt\ => \-stathalt\,
    stathenb => stathenb,
    \-step\ => \-step\,
    step => step,
    trapenb => trapenb
  );
  cadr_olord2_inst: cadr_olord2 port map (
      -- in ports
    aparok => aparok,
    \-busint.lm.reset\ => \-busint.lm.reset\,
    clk5 => clk5,
    dparok => dparok,
    errstop => errstop,
    \-halt\ => \-halt\,
    iparok => iparok,
    \-ldmode\ => \-ldmode\,
    mclk5 => mclk5,
    memparok => memparok,
    mmemparok => mmemparok,
    pdlparok => pdlparok,
    spcparok => spcparok,
    spy6 => spy6,
    spy7 => spy7,
    srun => srun,
    \stat.ovf\ => \stat.ovf\,
    \-upperhighok\ => \-upperhighok\,
    v0parok => v0parok,
    vmoparok => vmoparok,
      -- inout ports
    \-boot1\ => \-boot1\,
      -- out ports
    \-ape\ => \-ape\,
    \-boot\ => \-boot\,
    \boot.trap\ => \boot.trap\,
    \-boot2\ => \-boot2\,
    \bus.power.reset l\ => \bus.power.reset l\,
    \-bus.reset\ => \-bus.reset\,
    \-clk5\ => \-clk5\,
    clk5a => clk5a,
    \-clock reset a\ => \-clock reset a\,
    \-clock reset b\ => \-clock reset b\,
    \-dpe\ => \-dpe\,
    err => err,
    \-errhalt\ => \-errhalt\,
    \-halted\ => \-halted\,
    hi1 => hi1,
    hi2 => hi2,
    \-higherr\ => \-higherr\,
    highok => highok,
    \-ipe\ => \-ipe\,
    ldmode => ldmode,
    \-lowerhighok\ => \-lowerhighok\,
    \-mclk5\ => \-mclk5\,
    mclk5a => mclk5a,
    \-mempe\ => \-mempe\,
    \-mpe\ => \-mpe\,
    \-pdlpe\ => \-pdlpe\,
    \-power reset\ => \-power reset\,
    \power reset a\ => \power reset a\,
    \prog.boot\ => \prog.boot\,
    \prog.bus.reset\ => \prog.bus.reset\,
    \-prog.reset\ => \-prog.reset\,
    \-reset\ => \-reset\,
    reset => reset,
    \-spe\ => \-spe\,
    statstop => statstop,
    \-v0pe\ => \-v0pe\,
    \-v1pe\ => \-v1pe\
  );
  cadr_opcd_inst: cadr_opcd port map (
      -- in ports
    dc0 => dc0,
    dc1 => dc1,
    dc2 => dc2,
    dc3 => dc3,
    dc4 => dc4,
    dc5 => dc5,
    dc6 => dc6,
    dc7 => dc7,
    dc8 => dc8,
    dc9 => dc9,
    opc0 => opc0,
    opc1 => opc1,
    opc2 => opc2,
    opc3 => opc3,
    opc4 => opc4,
    opc5 => opc5,
    opc6 => opc6,
    opc7 => opc7,
    opc8 => opc8,
    opc9 => opc9,
    opc10 => opc10,
    opc11 => opc11,
    opc12 => opc12,
    opc13 => opc13,
    \-srcdc\ => \-srcdc\,
    \-srcopc\ => \-srcopc\,
    \-srcpdlidx\ => \-srcpdlidx\,
    \-srcpdlptr\ => \-srcpdlptr\,
    tse1b => tse1b,
      -- out ports
    dcdrive => dcdrive,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    \-opcdrive\ => \-opcdrive\,
    zero16 => zero16,
    \zero12.drive\ => \zero12.drive\,
    \-zero16.drive\ => \-zero16.drive\,
    \zero16.drive\ => \zero16.drive\
  );
  cadr_opcs_inst: cadr_opcs port map (
      -- in ports
    \-clk5\ => \-clk5\,
    hi2 => hi2,
    opcclk => opcclk,
    \-opcinh\ => \-opcinh\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
      -- out ports
    opc0 => opc0,
    opc1 => opc1,
    opc2 => opc2,
    opc3 => opc3,
    opc4 => opc4,
    opc5 => opc5,
    opc6 => opc6,
    opc7 => opc7,
    opc8 => opc8,
    opc9 => opc9,
    opc10 => opc10,
    opc11 => opc11,
    opc12 => opc12,
    opc13 => opc13,
    opcclka => opcclka,
    opcclkb => opcclkb,
    opcclkc => opcclkc,
    opcinha => opcinha,
    opcinhb => opcinhb
  );
  cadr_pctl_inst: cadr_pctl port map (
      -- in ports
    \-ape\ => \-ape\,
    \-dpe\ => \-dpe\,
    hi2 => hi2,
    \-idebug\ => \-idebug\,
    \-ipe\ => \-ipe\,
    \-iwriteda\ => \-iwriteda\,
    \-mempe\ => \-mempe\,
    \-mpe\ => \-mpe\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    \-pdlpe\ => \-pdlpe\,
    \-promdisabled\ => \-promdisabled\,
    \-spe\ => \-spe\,
    \-v0pe\ => \-v0pe\,
    \-v1pe\ => \-v1pe\,
      -- out ports
    \bottom.1k\ => \bottom.1k\,
    dpe => dpe,
    i46 => i46,
    ipe => ipe,
    \-promce0\ => \-promce0\,
    \-promce1\ => \-promce1\,
    \-promenable\ => \-promenable\,
    promenable => promenable,
    \-prompc0\ => \-prompc0\,
    \-prompc1\ => \-prompc1\,
    \-prompc2\ => \-prompc2\,
    \-prompc3\ => \-prompc3\,
    \-prompc4\ => \-prompc4\,
    \-prompc5\ => \-prompc5\,
    \-prompc6\ => \-prompc6\,
    \-prompc7\ => \-prompc7\,
    \-prompc8\ => \-prompc8\,
    \-prompc9\ => \-prompc9\,
    tilt0 => tilt0,
    tilt1 => tilt1
  );
  cadr_pdl0_inst: cadr_pdl0 port map (
      -- in ports
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
    \-pdla0b\ => \-pdla0b\,
    \-pdla1b\ => \-pdla1b\,
    \-pdla2b\ => \-pdla2b\,
    \-pdla3b\ => \-pdla3b\,
    \-pdla4b\ => \-pdla4b\,
    \-pdla5b\ => \-pdla5b\,
    \-pdla6b\ => \-pdla6b\,
    \-pdla7b\ => \-pdla7b\,
    \-pdla8b\ => \-pdla8b\,
    \-pdla9b\ => \-pdla9b\,
    \-pwpa\ => \-pwpa\,
    \-pwpb\ => \-pwpb\,
      -- out ports
    pdl16 => pdl16,
    pdl17 => pdl17,
    pdl18 => pdl18,
    pdl19 => pdl19,
    pdl20 => pdl20,
    pdl21 => pdl21,
    pdl22 => pdl22,
    pdl23 => pdl23,
    pdl24 => pdl24,
    pdl25 => pdl25,
    pdl26 => pdl26,
    pdl27 => pdl27,
    pdl28 => pdl28,
    pdl29 => pdl29,
    pdl30 => pdl30,
    pdl31 => pdl31,
    pdlparity => pdlparity
  );
  cadr_pdl1_inst: cadr_pdl1 port map (
      -- in ports
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    \-pdla0a\ => \-pdla0a\,
    \-pdla1a\ => \-pdla1a\,
    \-pdla2a\ => \-pdla2a\,
    \-pdla3a\ => \-pdla3a\,
    \-pdla4a\ => \-pdla4a\,
    \-pdla5a\ => \-pdla5a\,
    \-pdla6a\ => \-pdla6a\,
    \-pdla7a\ => \-pdla7a\,
    \-pdla8a\ => \-pdla8a\,
    \-pdla9a\ => \-pdla9a\,
    \-pwpb\ => \-pwpb\,
    \-pwpc\ => \-pwpc\,
      -- out ports
    pdl0 => pdl0,
    pdl1 => pdl1,
    pdl2 => pdl2,
    pdl3 => pdl3,
    pdl4 => pdl4,
    pdl5 => pdl5,
    pdl6 => pdl6,
    pdl7 => pdl7,
    pdl8 => pdl8,
    pdl9 => pdl9,
    pdl10 => pdl10,
    pdl11 => pdl11,
    pdl12 => pdl12,
    pdl13 => pdl13,
    pdl14 => pdl14,
    pdl15 => pdl15
  );
  cadr_pdlctl_inst: cadr_pdlctl port map (
      -- in ports
    clk4b => clk4b,
    \-clk4e\ => \-clk4e\,
    clk4f => clk4f,
    \-destpdl(p)\ => \-destpdl(p)\,
    \-destpdl(x)\ => \-destpdl(x)\,
    \-destpdltop\ => \-destpdltop\,
    \-destspc\ => \-destspc\,
    imod => imod,
    ir30 => ir30,
    nop => nop,
    pdlidx0 => pdlidx0,
    pdlidx1 => pdlidx1,
    pdlidx2 => pdlidx2,
    pdlidx3 => pdlidx3,
    pdlidx4 => pdlidx4,
    pdlidx5 => pdlidx5,
    pdlidx6 => pdlidx6,
    pdlidx7 => pdlidx7,
    pdlidx8 => pdlidx8,
    pdlidx9 => pdlidx9,
    pdlptr0 => pdlptr0,
    pdlptr1 => pdlptr1,
    pdlptr2 => pdlptr2,
    pdlptr3 => pdlptr3,
    pdlptr4 => pdlptr4,
    pdlptr5 => pdlptr5,
    pdlptr6 => pdlptr6,
    pdlptr7 => pdlptr7,
    pdlptr8 => pdlptr8,
    pdlptr9 => pdlptr9,
    \-reset\ => \-reset\,
    \-srcpdlpop\ => \-srcpdlpop\,
    \-srcpdltop\ => \-srcpdltop\,
    tse4b => tse4b,
    wp4a => wp4a,
      -- out ports
    \-destspcd\ => \-destspcd\,
    \-imodd\ => \-imodd\,
    imodd => imodd,
    \-pdla0a\ => \-pdla0a\,
    \-pdla0b\ => \-pdla0b\,
    \-pdla1a\ => \-pdla1a\,
    \-pdla1b\ => \-pdla1b\,
    \-pdla2a\ => \-pdla2a\,
    \-pdla2b\ => \-pdla2b\,
    \-pdla3a\ => \-pdla3a\,
    \-pdla3b\ => \-pdla3b\,
    \-pdla4a\ => \-pdla4a\,
    \-pdla4b\ => \-pdla4b\,
    \-pdla5a\ => \-pdla5a\,
    \-pdla5b\ => \-pdla5b\,
    \-pdla6a\ => \-pdla6a\,
    \-pdla6b\ => \-pdla6b\,
    \-pdla7a\ => \-pdla7a\,
    \-pdla7b\ => \-pdla7b\,
    \-pdla8a\ => \-pdla8a\,
    \-pdla8b\ => \-pdla8b\,
    \-pdla9a\ => \-pdla9a\,
    \-pdla9b\ => \-pdla9b\,
    \-pdlcnt\ => \-pdlcnt\,
    \-pdldrive\ => \-pdldrive\,
    pdlenb => pdlenb,
    \-pdlpa\ => \-pdlpa\,
    \-pdlpb\ => \-pdlpb\,
    pdlwrite => pdlwrite,
    \-pdlwrited\ => \-pdlwrited\,
    pdlwrited => pdlwrited,
    \-pwidx\ => \-pwidx\,
    pwidx => pwidx,
    \-pwpa\ => \-pwpa\,
    \-pwpb\ => \-pwpb\,
    \-pwpc\ => \-pwpc\
  );
  cadr_pdlptr_inst: cadr_pdlptr port map (
      -- in ports
    clk3f => clk3f,
    \-destpdlp\ => \-destpdlp\,
    \-destpdlx\ => \-destpdlx\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    \-pdlcnt\ => \-pdlcnt\,
    srcpdlidx => srcpdlidx,
    \-srcpdlpop\ => \-srcpdlpop\,
    srcpdlptr => srcpdlptr,
    tse4b => tse4b,
      -- out ports
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    \-pdlcry3\ => \-pdlcry3\,
    \-pdlcry7\ => \-pdlcry7\,
    pdlidx0 => pdlidx0,
    pdlidx1 => pdlidx1,
    pdlidx2 => pdlidx2,
    pdlidx3 => pdlidx3,
    pdlidx4 => pdlidx4,
    pdlidx5 => pdlidx5,
    pdlidx6 => pdlidx6,
    pdlidx7 => pdlidx7,
    pdlidx8 => pdlidx8,
    pdlidx9 => pdlidx9,
    pdlptr0 => pdlptr0,
    pdlptr1 => pdlptr1,
    pdlptr2 => pdlptr2,
    pdlptr3 => pdlptr3,
    pdlptr4 => pdlptr4,
    pdlptr5 => pdlptr5,
    pdlptr6 => pdlptr6,
    pdlptr7 => pdlptr7,
    pdlptr8 => pdlptr8,
    pdlptr9 => pdlptr9,
    pidrive => pidrive,
    \-ppdrive\ => \-ppdrive\
  );
  cadr_platch_inst: cadr_platch port map (
      -- in ports
    clk4a => clk4a,
    pdl0 => pdl0,
    pdl1 => pdl1,
    pdl2 => pdl2,
    pdl3 => pdl3,
    pdl4 => pdl4,
    pdl5 => pdl5,
    pdl6 => pdl6,
    pdl7 => pdl7,
    pdl8 => pdl8,
    pdl9 => pdl9,
    pdl10 => pdl10,
    pdl11 => pdl11,
    pdl12 => pdl12,
    pdl13 => pdl13,
    pdl14 => pdl14,
    pdl15 => pdl15,
    pdl16 => pdl16,
    pdl17 => pdl17,
    pdl18 => pdl18,
    pdl19 => pdl19,
    pdl20 => pdl20,
    pdl21 => pdl21,
    pdl22 => pdl22,
    pdl23 => pdl23,
    pdl24 => pdl24,
    pdl25 => pdl25,
    pdl26 => pdl26,
    pdl27 => pdl27,
    pdl28 => pdl28,
    pdl29 => pdl29,
    pdl30 => pdl30,
    pdl31 => pdl31,
    \-pdldrive\ => \-pdldrive\,
    pdlparity => pdlparity,
      -- out ports
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    mparity => mparity
  );
  cadr_prom0_inst: cadr_prom0 port map (
      -- in ports
    \-promce0\ => \-promce0\,
    \-prompc0\ => \-prompc0\,
    \-prompc1\ => \-prompc1\,
    \-prompc2\ => \-prompc2\,
    \-prompc3\ => \-prompc3\,
    \-prompc4\ => \-prompc4\,
    \-prompc5\ => \-prompc5\,
    \-prompc6\ => \-prompc6\,
    \-prompc7\ => \-prompc7\,
    \-prompc8\ => \-prompc8\,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i47 => i47,
    i48 => i48
  );
  cadr_prom1_inst: cadr_prom1 port map (
      -- in ports
    \-promce1\ => \-promce1\,
    \-prompc0\ => \-prompc0\,
    \-prompc1\ => \-prompc1\,
    \-prompc2\ => \-prompc2\,
    \-prompc3\ => \-prompc3\,
    \-prompc4\ => \-prompc4\,
    \-prompc5\ => \-prompc5\,
    \-prompc6\ => \-prompc6\,
    \-prompc7\ => \-prompc7\,
    \-prompc8\ => \-prompc8\,
      -- out ports
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i47 => i47,
    i48 => i48
  );
  cadr_q_inst: cadr_q port map (
      -- in ports
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    \-alu31\ => \-alu31\,
    alu31 => alu31,
    clk2b => clk2b,
    hi7 => hi7,
    qs0 => qs0,
    qs1 => qs1,
      -- out ports
    q0 => q0,
    q1 => q1,
    q2 => q2,
    q3 => q3,
    q4 => q4,
    q5 => q5,
    q6 => q6,
    q7 => q7,
    q8 => q8,
    q9 => q9,
    q10 => q10,
    q11 => q11,
    q12 => q12,
    q13 => q13,
    q14 => q14,
    q15 => q15,
    q16 => q16,
    q17 => q17,
    q18 => q18,
    q19 => q19,
    q20 => q20,
    q21 => q21,
    q22 => q22,
    q23 => q23,
    q24 => q24,
    q25 => q25,
    q26 => q26,
    q27 => q27,
    q28 => q28,
    q29 => q29,
    q30 => q30,
    q31 => q31
  );
  cadr_qctl_inst: cadr_qctl port map (
      -- in ports
    alu31 => alu31,
    \-ir0\ => \-ir0\,
    \-ir1\ => \-ir1\,
    \-iralu\ => \-iralu\,
    q0 => q0,
    q1 => q1,
    q2 => q2,
    q3 => q3,
    q4 => q4,
    q5 => q5,
    q6 => q6,
    q7 => q7,
    q8 => q8,
    q9 => q9,
    q10 => q10,
    q11 => q11,
    q12 => q12,
    q13 => q13,
    q14 => q14,
    q15 => q15,
    q16 => q16,
    q17 => q17,
    q18 => q18,
    q19 => q19,
    q20 => q20,
    q21 => q21,
    q22 => q22,
    q23 => q23,
    q24 => q24,
    q25 => q25,
    q26 => q26,
    q27 => q27,
    q28 => q28,
    q29 => q29,
    q30 => q30,
    q31 => q31,
    \-srcq\ => \-srcq\,
    tse2 => tse2,
      -- out ports
    \-alu31\ => \-alu31\,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    \-qdrive\ => \-qdrive\,
    qdrive => qdrive,
    qs0 => qs0,
    qs1 => qs1,
    srcq => srcq
  );
  cadr_shift0_inst: cadr_shift0 port map (
      -- in ports
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    s0 => s0,
    s1 => s1,
    \-s4\ => \-s4\,
    s4 => s4,
    s2a => s2a,
    s3a => s3a,
    sa16 => sa16,
    sa17 => sa17,
    sa18 => sa18,
    sa19 => sa19,
    sa20 => sa20,
    sa21 => sa21,
    sa22 => sa22,
    sa23 => sa23,
    sa24 => sa24,
    sa25 => sa25,
    sa26 => sa26,
    sa27 => sa27,
    sa28 => sa28,
    sa29 => sa29,
    sa30 => sa30,
    sa31 => sa31,
      -- out ports
    m5 => m5,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    r7 => r7,
    r8 => r8,
    r9 => r9,
    r10 => r10,
    r11 => r11,
    r12 => r12,
    r13 => r13,
    r14 => r14,
    r15 => r15,
    sa0 => sa0,
    sa1 => sa1,
    sa2 => sa2,
    sa3 => sa3,
    sa4 => sa4,
    sa5 => sa5,
    sa6 => sa6,
    sa7 => sa7,
    sa8 => sa8,
    sa9 => sa9,
    sa10 => sa10,
    sa11 => sa11,
    sa12 => sa12,
    sa13 => sa13,
    sa14 => sa14,
    sa15 => sa15
  );
  cadr_shift1_inst: cadr_shift1 port map (
      -- in ports
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    s0 => s0,
    s1 => s1,
    \-s4\ => \-s4\,
    s4 => s4,
    s2b => s2b,
    s3b => s3b,
    sa0 => sa0,
    sa1 => sa1,
    sa2 => sa2,
    sa3 => sa3,
    sa4 => sa4,
    sa5 => sa5,
    sa6 => sa6,
    sa7 => sa7,
    sa8 => sa8,
    sa9 => sa9,
    sa10 => sa10,
    sa11 => sa11,
    sa12 => sa12,
    sa13 => sa13,
    sa14 => sa14,
    sa15 => sa15,
      -- out ports
    r16 => r16,
    r17 => r17,
    r18 => r18,
    r19 => r19,
    r20 => r20,
    r21 => r21,
    r22 => r22,
    r23 => r23,
    r24 => r24,
    r25 => r25,
    r26 => r26,
    r27 => r27,
    r28 => r28,
    r29 => r29,
    r30 => r30,
    r31 => r31,
    sa16 => sa16,
    sa17 => sa17,
    sa18 => sa18,
    sa19 => sa19,
    sa20 => sa20,
    sa21 => sa21,
    sa22 => sa22,
    sa23 => sa23,
    sa24 => sa24,
    sa25 => sa25,
    sa26 => sa26,
    sa27 => sa27,
    sa28 => sa28,
    sa29 => sa29,
    sa30 => sa30,
    sa31 => sa31
  );
  cadr_smctl_inst: cadr_smctl port map (
      -- in ports
    \-ir0\ => \-ir0\,
    \-ir1\ => \-ir1\,
    \-ir2\ => \-ir2\,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir12 => ir12,
    ir13 => ir13,
    \-irbyte\ => \-irbyte\,
    \-sh3\ => \-sh3\,
    \-sh4\ => \-sh4\,
      -- out ports
    \-mr\ => \-mr\,
    mskl0 => mskl0,
    mskl1 => mskl1,
    mskl2 => mskl2,
    mskl3 => mskl3,
    mskl4 => mskl4,
    mskl3cry => mskl3cry,
    mskr0 => mskr0,
    mskr1 => mskr1,
    mskr2 => mskr2,
    mskr3 => mskr3,
    mskr4 => mskr4,
    s0 => s0,
    s1 => s1,
    \-s4\ => \-s4\,
    s4 => s4,
    s2a => s2a,
    s2b => s2b,
    s3a => s3a,
    s3b => s3b,
    \-sr\ => \-sr\
  );
  cadr_source_inst: cadr_source port map (
      -- in ports
    hi5 => hi5,
    \-idebug\ => \-idebug\,
    ir3 => ir3,
    ir4 => ir4,
    ir8 => ir8,
    ir10 => ir10,
    ir11 => ir11,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    \-ir31\ => \-ir31\,
    ir43 => ir43,
    ir44 => ir44,
    \-iwrited\ => \-iwrited\,
    nop => nop,
      -- out ports
    dest => dest,
    \-destimod0\ => \-destimod0\,
    \-destimod1\ => \-destimod1\,
    \-destintctl\ => \-destintctl\,
    \-destlc\ => \-destlc\,
    destm => destm,
    \-destmdr\ => \-destmdr\,
    \-destmem\ => \-destmem\,
    \-destpdl(p)\ => \-destpdl(p)\,
    \-destpdl(x)\ => \-destpdl(x)\,
    \-destpdlp\ => \-destpdlp\,
    \-destpdltop\ => \-destpdltop\,
    \-destpdlx\ => \-destpdlx\,
    \-destspc\ => \-destspc\,
    \-destvma\ => \-destvma\,
    \-div\ => \-div\,
    \-funct0\ => \-funct0\,
    \-funct1\ => \-funct1\,
    \-funct2\ => \-funct2\,
    \-funct3\ => \-funct3\,
    imod => imod,
    \-ir22\ => \-ir22\,
    \-ir25\ => \-ir25\,
    \-iralu\ => \-iralu\,
    iralu => iralu,
    \-irbyte\ => \-irbyte\,
    \-irdisp\ => \-irdisp\,
    irdisp => irdisp,
    \-irjump\ => \-irjump\,
    irjump => irjump,
    \-mul\ => \-mul\,
    \-specalu\ => \-specalu\,
    \-srcdc\ => \-srcdc\,
    \-srclc\ => \-srclc\,
    \-srcmap\ => \-srcmap\,
    \-srcmd\ => \-srcmd\,
    \-srcopc\ => \-srcopc\,
    \-srcpdlidx\ => \-srcpdlidx\,
    \-srcpdlpop\ => \-srcpdlpop\,
    \-srcpdlptr\ => \-srcpdlptr\,
    \-srcpdltop\ => \-srcpdltop\,
    \-srcq\ => \-srcq\,
    \-srcspc\ => \-srcspc\,
    \-srcspcpop\ => \-srcspcpop\,
    \-srcvma\ => \-srcvma\
  );
  cadr_spc_inst: cadr_spc port map (
      -- in ports
    clk4f => clk4f,
    \-spcnt\ => \-spcnt\,
    spcw0 => spcw0,
    spcw1 => spcw1,
    spcw2 => spcw2,
    spcw3 => spcw3,
    spcw4 => spcw4,
    spcw5 => spcw5,
    spcw6 => spcw6,
    spcw7 => spcw7,
    spcw8 => spcw8,
    spcw9 => spcw9,
    spcw10 => spcw10,
    spcw11 => spcw11,
    spcw12 => spcw12,
    spcw13 => spcw13,
    spcw14 => spcw14,
    spcw15 => spcw15,
    spcw16 => spcw16,
    spcw17 => spcw17,
    spcw18 => spcw18,
    spcwpar => spcwpar,
    spush => spush,
    \-swpa\ => \-swpa\,
    \-swpb\ => \-swpb\,
      -- out ports
    hi1 => hi1,
    hi2 => hi2,
    hi3 => hi3,
    hi4 => hi4,
    hi5 => hi5,
    hi6 => hi6,
    hi7 => hi7,
    hi8 => hi8,
    hi9 => hi9,
    hi10 => hi10,
    hi11 => hi11,
    hi12 => hi12,
    \-spccry\ => \-spccry\,
    spco0 => spco0,
    spco1 => spco1,
    spco2 => spco2,
    spco3 => spco3,
    spco4 => spco4,
    spco5 => spco5,
    spco6 => spco6,
    spco7 => spco7,
    spco8 => spco8,
    spco9 => spco9,
    spco10 => spco10,
    spco11 => spco11,
    spco12 => spco12,
    spco13 => spco13,
    spco14 => spco14,
    spco15 => spco15,
    spco16 => spco16,
    spco17 => spco17,
    spco18 => spco18,
    spcopar => spcopar,
    spcptr0 => spcptr0,
    spcptr1 => spcptr1,
    spcptr2 => spcptr2,
    spcptr3 => spcptr3,
    spcptr4 => spcptr4
  );
  cadr_spclch_inst: cadr_spclch port map (
      -- in ports
    clk4c => clk4c,
    clk4d => clk4d,
    hi1 => hi1,
    \-spcdrive\ => \-spcdrive\,
    spcdrive => spcdrive,
    spco0 => spco0,
    spco1 => spco1,
    spco2 => spco2,
    spco3 => spco3,
    spco4 => spco4,
    spco5 => spco5,
    spco6 => spco6,
    spco7 => spco7,
    spco8 => spco8,
    spco9 => spco9,
    spco10 => spco10,
    spco11 => spco11,
    spco12 => spco12,
    spco13 => spco13,
    spco14 => spco14,
    spco15 => spco15,
    spco16 => spco16,
    spco17 => spco17,
    spco18 => spco18,
    spcopar => spcopar,
    \-spcpass\ => \-spcpass\,
    spcptr0 => spcptr0,
    spcptr1 => spcptr1,
    spcptr2 => spcptr2,
    spcptr3 => spcptr3,
    spcptr4 => spcptr4,
    spcw0 => spcw0,
    spcw1 => spcw1,
    spcw2 => spcw2,
    spcw3 => spcw3,
    spcw4 => spcw4,
    spcw5 => spcw5,
    spcw6 => spcw6,
    spcw7 => spcw7,
    spcw8 => spcw8,
    spcw9 => spcw9,
    spcw10 => spcw10,
    spcw11 => spcw11,
    spcw12 => spcw12,
    spcw13 => spcw13,
    spcw14 => spcw14,
    spcw15 => spcw15,
    spcw16 => spcw16,
    spcw17 => spcw17,
    spcw18 => spcw18,
    spcwpar => spcwpar,
    \-spcwpass\ => \-spcwpass\,
    spcwpass => spcwpass,
      -- out ports
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    spc0 => spc0,
    spc1 => spc1,
    spc2 => spc2,
    spc3 => spc3,
    spc4 => spc4,
    spc5 => spc5,
    spc6 => spc6,
    spc7 => spc7,
    spc8 => spc8,
    spc9 => spc9,
    spc10 => spc10,
    spc11 => spc11,
    spc12 => spc12,
    spc13 => spc13,
    spc14 => spc14,
    spc15 => spc15,
    spc16 => spc16,
    spc17 => spc17,
    spc18 => spc18,
    spcpar => spcpar
  );
  cadr_spcpar_inst: cadr_spcpar port map (
      -- in ports
    spc0 => spc0,
    spc1 => spc1,
    spc2 => spc2,
    spc3 => spc3,
    spc4 => spc4,
    spc5 => spc5,
    spc6 => spc6,
    spc7 => spc7,
    spc8 => spc8,
    spc9 => spc9,
    spc10 => spc10,
    spc11 => spc11,
    spc12 => spc12,
    spc13 => spc13,
    spc14 => spc14,
    spc15 => spc15,
    spc16 => spc16,
    spc17 => spc17,
    spc18 => spc18,
    spcpar => spcpar,
    spcw0 => spcw0,
    spcw1 => spcw1,
    spcw2 => spcw2,
    spcw3 => spcw3,
    spcw4 => spcw4,
    spcw5 => spcw5,
    spcw6 => spcw6,
    spcw7 => spcw7,
    spcw8 => spcw8,
    spcw9 => spcw9,
    spcw10 => spcw10,
    spcw11 => spcw11,
    spcw12 => spcw12,
    spcw13 => spcw13,
    spcw14 => spcw14,
    spcw15 => spcw15,
    spcw16 => spcw16,
    spcw17 => spcw17,
    spcw18 => spcw18,
      -- out ports
    spcparh => spcparh,
    spcparok => spcparok,
    spcwpar => spcwpar,
    spcwparh => spcwparh,
    \-spcwparl\ => \-spcwparl\
  );
  cadr_spcw_inst: cadr_spcw port map (
      -- in ports
    clk4d => clk4d,
    destspcd => destspcd,
    ipc0 => ipc0,
    ipc1 => ipc1,
    ipc2 => ipc2,
    ipc3 => ipc3,
    ipc4 => ipc4,
    ipc5 => ipc5,
    ipc6 => ipc6,
    ipc7 => ipc7,
    ipc8 => ipc8,
    ipc9 => ipc9,
    ipc10 => ipc10,
    ipc11 => ipc11,
    ipc12 => ipc12,
    ipc13 => ipc13,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    n => n,
    wpc0 => wpc0,
    wpc1 => wpc1,
    wpc2 => wpc2,
    wpc3 => wpc3,
    wpc4 => wpc4,
    wpc5 => wpc5,
    wpc6 => wpc6,
    wpc7 => wpc7,
    wpc8 => wpc8,
    wpc9 => wpc9,
    wpc10 => wpc10,
    wpc11 => wpc11,
    wpc12 => wpc12,
    wpc13 => wpc13,
      -- out ports
    reta0 => reta0,
    reta1 => reta1,
    reta2 => reta2,
    reta3 => reta3,
    reta4 => reta4,
    reta5 => reta5,
    reta6 => reta6,
    reta7 => reta7,
    reta8 => reta8,
    reta9 => reta9,
    reta10 => reta10,
    reta11 => reta11,
    reta12 => reta12,
    reta13 => reta13,
    spcw0 => spcw0,
    spcw1 => spcw1,
    spcw2 => spcw2,
    spcw3 => spcw3,
    spcw4 => spcw4,
    spcw5 => spcw5,
    spcw6 => spcw6,
    spcw7 => spcw7,
    spcw8 => spcw8,
    spcw9 => spcw9,
    spcw10 => spcw10,
    spcw11 => spcw11,
    spcw12 => spcw12,
    spcw13 => spcw13,
    spcw14 => spcw14,
    spcw15 => spcw15,
    spcw16 => spcw16,
    spcw17 => spcw17,
    spcw18 => spcw18
  );
  cadr_spy0_inst: cadr_spy0 port map (
      -- in ports
    \-dbread\ => \-dbread\,
    \-dbwrite\ => \-dbwrite\,
    eadr0 => eadr0,
    eadr1 => eadr1,
    eadr2 => eadr2,
    eadr3 => eadr3,
    hi1 => hi1,
      -- out ports
    \-ldclk\ => \-ldclk\,
    \-lddbirh\ => \-lddbirh\,
    \-lddbirl\ => \-lddbirl\,
    \-lddbirm\ => \-lddbirm\,
    \-ldmode\ => \-ldmode\,
    \-ldopc\ => \-ldopc\,
    \-spy.ah\ => \-spy.ah\,
    \-spy.al\ => \-spy.al\,
    \-spy.flag1\ => \-spy.flag1\,
    \-spy.flag2\ => \-spy.flag2\,
    \-spy.irh\ => \-spy.irh\,
    \-spy.irl\ => \-spy.irl\,
    \-spy.irm\ => \-spy.irm\,
    \-spy.mh\ => \-spy.mh\,
    \-spy.ml\ => \-spy.ml\,
    \-spy.obh\ => \-spy.obh\,
    \-spy.obl\ => \-spy.obl\,
    \-spy.opc\ => \-spy.opc\,
    \-spy.pc\ => \-spy.pc\,
    \-spy.sth\ => \-spy.sth\,
    \-spy.stl\ => \-spy.stl\
  );
  cadr_spy1_inst: cadr_spy1 port map (
      -- in ports
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir10 => ir10,
    ir11 => ir11,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    ir31 => ir31,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    ir42 => ir42,
    ir43 => ir43,
    ir44 => ir44,
    ir45 => ir45,
    ir46 => ir46,
    ir47 => ir47,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    \-spy.irh\ => \-spy.irh\,
    \-spy.irl\ => \-spy.irl\,
    \-spy.irm\ => \-spy.irm\,
    \-spy.obh\ => \-spy.obh\,
      -- out ports
    \-spy.obl\ => \-spy.obl\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15
  );
  cadr_spy2_inst: cadr_spy2 port map (
      -- in ports
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    destspcd => destspcd,
    imodd => imodd,
    ir48 => ir48,
    iwrited => iwrited,
    jcond => jcond,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    nop => nop,
    pcs0 => pcs0,
    pcs1 => pcs1,
    pdlwrited => pdlwrited,
    spushd => spushd,
    \-spy.ah\ => \-spy.ah\,
    \-spy.flag2\ => \-spy.flag2\,
    \-spy.mh\ => \-spy.mh\,
    \-spy.ml\ => \-spy.ml\,
    \-vmaok\ => \-vmaok\,
    wmapd => wmapd,
      -- out ports
    \-spy.al\ => \-spy.al\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15
  );
  cadr_spy4_inst: cadr_spy4 port map (
      -- in ports
    \-ape\ => \-ape\,
    \-dpe\ => \-dpe\,
    err => err,
    \-higherr\ => \-higherr\,
    \-ipe\ => \-ipe\,
    \-mempe\ => \-mempe\,
    \-mpe\ => \-mpe\,
    opc0 => opc0,
    opc1 => opc1,
    opc2 => opc2,
    opc3 => opc3,
    opc4 => opc4,
    opc5 => opc5,
    opc6 => opc6,
    opc7 => opc7,
    opc8 => opc8,
    opc9 => opc9,
    opc10 => opc10,
    opc11 => opc11,
    opc12 => opc12,
    opc13 => opc13,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    \-pdlpe\ => \-pdlpe\,
    promdisable => promdisable,
    \-spe\ => \-spe\,
    \-spy.opc\ => \-spy.opc\,
    \-spy.pc\ => \-spy.pc\,
    srun => srun,
    ssdone => ssdone,
    \-stathalt\ => \-stathalt\,
    \-v0pe\ => \-v0pe\,
    \-v1pe\ => \-v1pe\,
    \-wait\ => \-wait\,
      -- out ports
    \-spy.flag1\ => \-spy.flag1\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15
  );
  cadr_stat_inst: cadr_stat port map (
      -- in ports
    clk5a => clk5a,
    hi1 => hi1,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    \-ldstat\ => \-ldstat\,
    \-spy.sth\ => \-spy.sth\,
    \-spy.stl\ => \-spy.stl\,
    \-statbit\ => \-statbit\,
      -- out ports
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15,
    st0 => st0,
    st1 => st1,
    st2 => st2,
    st3 => st3,
    st4 => st4,
    st5 => st5,
    st6 => st6,
    st7 => st7,
    st8 => st8,
    st9 => st9,
    st10 => st10,
    st11 => st11,
    st12 => st12,
    st13 => st13,
    st14 => st14,
    st15 => st15,
    st16 => st16,
    st17 => st17,
    st18 => st18,
    st19 => st19,
    st20 => st20,
    st21 => st21,
    st22 => st22,
    st23 => st23,
    st24 => st24,
    st25 => st25,
    st26 => st26,
    st27 => st27,
    st28 => st28,
    st29 => st29,
    st30 => st30,
    st31 => st31,
    \-stc4\ => \-stc4\,
    \-stc8\ => \-stc8\,
    \-stc12\ => \-stc12\,
    \-stc16\ => \-stc16\,
    \-stc20\ => \-stc20\,
    \-stc24\ => \-stc24\,
    \-stc28\ => \-stc28\,
    \-stc32\ => \-stc32\
  );
  cadr_trap_inst: cadr_trap port map (
      -- in ports
    \boot.trap\ => \boot.trap\,
    \-md0\ => \-md0\,
    \-md1\ => \-md1\,
    \-md2\ => \-md2\,
    \-md3\ => \-md3\,
    \-md4\ => \-md4\,
    \-md5\ => \-md5\,
    \-md6\ => \-md6\,
    \-md7\ => \-md7\,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-md24\ => \-md24\,
    \-md25\ => \-md25\,
    \-md26\ => \-md26\,
    \-md27\ => \-md27\,
    \-md28\ => \-md28\,
    \-md29\ => \-md29\,
    \-md30\ => \-md30\,
    \-md31\ => \-md31\,
    mdhaspar => mdhaspar,
    mdpar => mdpar,
    trapenb => trapenb,
    \use.md\ => \use.md\,
    \-wait\ => \-wait\,
      -- out ports
    mdparerr => mdparerr,
    mdpareven => mdpareven,
    mdparl => mdparl,
    mdparm => mdparm,
    mdparodd => mdparodd,
    \-memparok\ => \-memparok\,
    memparok => memparok,
    \-parerr\ => \-parerr\,
    \-trap\ => \-trap\,
    trapa => trapa,
    trapb => trapb,
    \-trapenb\ => \-trapenb\
  );
  cadr_vctl1_inst: cadr_vctl1 port map (
      -- in ports
    clk2a => clk2a,
    clk2c => clk2c,
    \-clk3g\ => \-clk3g\,
    destmem => destmem,
    hi4 => hi4,
    hi11 => hi11,
    \-ifetch\ => \-ifetch\,
    lcinc => lcinc,
    \-lvmo22\ => \-lvmo22\,
    mclk1a => mclk1a,
    \-memack\ => \-memack\,
    \-memgrant\ => \-memgrant\,
    \-memprepare\ => \-memprepare\,
    \-memrd\ => \-memrd\,
    \-memwr\ => \-memwr\,
    needfetch => needfetch,
    \-pfr\ => \-pfr\,
    \-reset\ => \-reset\,
    \use.md\ => \use.md\,
    wmap => wmap,
      -- out ports
    \-hang\ => \-hang\,
    mbusy => mbusy,
    \-mbusy.sync\ => \-mbusy.sync\,
    \mbusy.sync\ => \mbusy.sync\,
    \-memop\ => \-memop\,
    memprepare => memprepare,
    memrq => memrq,
    \-memstart\ => \-memstart\,
    memstart => memstart,
    \-mfinish\ => \-mfinish\,
    \-mfinishd\ => \-mfinishd\,
    \-pfw\ => \-pfw\,
    \rd.in.progress\ => \rd.in.progress\,
    rdcyc => rdcyc,
    \-rdfinish\ => \-rdfinish\,
    \set.rd.in.progress\ => \set.rd.in.progress\,
    \-vmaok\ => \-vmaok\,
    \-wait\ => \-wait\,
    \-wmapd\ => \-wmapd\,
    wmapd => wmapd,
    wrcyc => wrcyc
  );
  cadr_vctl2_inst: cadr_vctl2 port map (
      -- in ports
    clk2c => clk2c,
    \-destmdr\ => \-destmdr\,
    \-destmem\ => \-destmem\,
    \-destvma\ => \-destvma\,
    hi11 => hi11,
    \-ifetch\ => \-ifetch\,
    ir19 => ir19,
    ir20 => ir20,
    \lm drive enb\ => \lm drive enb\,
    \-lvmo23\ => \-lvmo23\,
    memprepare => memprepare,
    memrq => memrq,
    \-nopa\ => \-nopa\,
    \-srcmd\ => \-srcmd\,
    \-vma25\ => \-vma25\,
    \-vma26\ => \-vma26\,
    wp1a => wp1a,
    wp1b => wp1b,
    wrcyc => wrcyc,
      -- out ports
    destmem => destmem,
    mapwr0d => mapwr0d,
    mapwr1d => mapwr1d,
    mdsela => mdsela,
    mdselb => mdselb,
    \-memdrive.a\ => \-memdrive.a\,
    \-memdrive.b\ => \-memdrive.b\,
    \-memprepare\ => \-memprepare\,
    \-memrd\ => \-memrd\,
    \-memrq\ => \-memrq\,
    \-memwr\ => \-memwr\,
    nopa => nopa,
    \-pfr\ => \-pfr\,
    \use.md\ => \use.md\,
    \-vm0wpa\ => \-vm0wpa\,
    \-vm0wpb\ => \-vm0wpb\,
    \-vm1wpa\ => \-vm1wpa\,
    \-vm1wpb\ => \-vm1wpb\,
    \-vmaenb\ => \-vmaenb\,
    vmasela => vmasela,
    vmaselb => vmaselb,
    \-wmap\ => \-wmap\,
    wmap => wmap,
    \-wmapd\ => \-wmapd\
  );
  cadr_vma_inst: cadr_vma port map (
      -- in ports
    clk1a => clk1a,
    clk2a => clk2a,
    clk2c => clk2c,
    \-srcvma\ => \-srcvma\,
    tse2 => tse2,
    \-vmaenb\ => \-vmaenb\,
    \-vmas0\ => \-vmas0\,
    \-vmas1\ => \-vmas1\,
    \-vmas2\ => \-vmas2\,
    \-vmas3\ => \-vmas3\,
    \-vmas4\ => \-vmas4\,
    \-vmas5\ => \-vmas5\,
    \-vmas6\ => \-vmas6\,
    \-vmas7\ => \-vmas7\,
    \-vmas8\ => \-vmas8\,
    \-vmas9\ => \-vmas9\,
    \-vmas10\ => \-vmas10\,
    \-vmas11\ => \-vmas11\,
    \-vmas12\ => \-vmas12\,
    \-vmas13\ => \-vmas13\,
    \-vmas14\ => \-vmas14\,
    \-vmas15\ => \-vmas15\,
    \-vmas16\ => \-vmas16\,
    \-vmas17\ => \-vmas17\,
    \-vmas18\ => \-vmas18\,
    \-vmas19\ => \-vmas19\,
    \-vmas20\ => \-vmas20\,
    \-vmas21\ => \-vmas21\,
    \-vmas22\ => \-vmas22\,
    \-vmas23\ => \-vmas23\,
    \-vmas24\ => \-vmas24\,
    \-vmas25\ => \-vmas25\,
    \-vmas26\ => \-vmas26\,
    \-vmas27\ => \-vmas27\,
    \-vmas28\ => \-vmas28\,
    \-vmas29\ => \-vmas29\,
    \-vmas30\ => \-vmas30\,
    \-vmas31\ => \-vmas31\,
      -- out ports
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    srcvma => srcvma,
    \-vma0\ => \-vma0\,
    \-vma1\ => \-vma1\,
    \-vma2\ => \-vma2\,
    \-vma3\ => \-vma3\,
    \-vma4\ => \-vma4\,
    \-vma5\ => \-vma5\,
    \-vma6\ => \-vma6\,
    \-vma7\ => \-vma7\,
    \-vma8\ => \-vma8\,
    \-vma9\ => \-vma9\,
    \-vma10\ => \-vma10\,
    \-vma11\ => \-vma11\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    \-vma24\ => \-vma24\,
    \-vma25\ => \-vma25\,
    \-vma26\ => \-vma26\,
    \-vma27\ => \-vma27\,
    \-vma28\ => \-vma28\,
    \-vma29\ => \-vma29\,
    \-vma30\ => \-vma30\,
    \-vma31\ => \-vma31\,
    \-vmadrive\ => \-vmadrive\
  );
  cadr_vmas_inst: cadr_vmas port map (
      -- in ports
    lc2 => lc2,
    lc3 => lc3,
    lc4 => lc4,
    lc5 => lc5,
    lc6 => lc6,
    lc7 => lc7,
    lc8 => lc8,
    lc9 => lc9,
    lc10 => lc10,
    lc11 => lc11,
    lc12 => lc12,
    lc13 => lc13,
    lc14 => lc14,
    lc15 => lc15,
    lc16 => lc16,
    lc17 => lc17,
    lc18 => lc18,
    lc19 => lc19,
    lc20 => lc20,
    lc21 => lc21,
    lc22 => lc22,
    lc23 => lc23,
    lc24 => lc24,
    lc25 => lc25,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-memstart\ => \-memstart\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    \-vma8\ => \-vma8\,
    \-vma9\ => \-vma9\,
    \-vma10\ => \-vma10\,
    \-vma11\ => \-vma11\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    vmasela => vmasela,
    vmaselb => vmaselb,
      -- out ports
    mapi8 => mapi8,
    mapi9 => mapi9,
    mapi10 => mapi10,
    mapi11 => mapi11,
    mapi12 => mapi12,
    mapi13 => mapi13,
    mapi14 => mapi14,
    mapi15 => mapi15,
    mapi16 => mapi16,
    mapi17 => mapi17,
    mapi18 => mapi18,
    mapi19 => mapi19,
    mapi20 => mapi20,
    mapi21 => mapi21,
    mapi22 => mapi22,
    mapi23 => mapi23,
    \-vmas0\ => \-vmas0\,
    \-vmas1\ => \-vmas1\,
    \-vmas2\ => \-vmas2\,
    \-vmas3\ => \-vmas3\,
    \-vmas4\ => \-vmas4\,
    \-vmas5\ => \-vmas5\,
    \-vmas6\ => \-vmas6\,
    \-vmas7\ => \-vmas7\,
    \-vmas8\ => \-vmas8\,
    \-vmas9\ => \-vmas9\,
    \-vmas10\ => \-vmas10\,
    \-vmas11\ => \-vmas11\,
    \-vmas12\ => \-vmas12\,
    \-vmas13\ => \-vmas13\,
    \-vmas14\ => \-vmas14\,
    \-vmas15\ => \-vmas15\,
    \-vmas16\ => \-vmas16\,
    \-vmas17\ => \-vmas17\,
    \-vmas18\ => \-vmas18\,
    \-vmas19\ => \-vmas19\,
    \-vmas20\ => \-vmas20\,
    \-vmas21\ => \-vmas21\,
    \-vmas22\ => \-vmas22\,
    \-vmas23\ => \-vmas23\,
    \-vmas24\ => \-vmas24\,
    \-vmas25\ => \-vmas25\,
    \-vmas26\ => \-vmas26\,
    \-vmas27\ => \-vmas27\,
    \-vmas28\ => \-vmas28\,
    \-vmas29\ => \-vmas29\,
    \-vmas30\ => \-vmas30\,
    \-vmas31\ => \-vmas31\
  );
  cadr_vmem0_inst: cadr_vmem0 port map (
      -- in ports
    mapi13 => mapi13,
    mapi14 => mapi14,
    mapi15 => mapi15,
    mapi16 => mapi16,
    mapi17 => mapi17,
    mapi18 => mapi18,
    mapi19 => mapi19,
    mapi20 => mapi20,
    mapi21 => mapi21,
    mapi22 => mapi22,
    mapi23 => mapi23,
    memstart => memstart,
    srcmap => srcmap,
    \-vm0wpa\ => \-vm0wpa\,
    \-vm0wpb\ => \-vm0wpb\,
    \-vma27\ => \-vma27\,
    \-vma28\ => \-vma28\,
    \-vma29\ => \-vma29\,
    \-vma30\ => \-vma30\,
    \-vma31\ => \-vma31\,
    vmoparodd => vmoparodd,
      -- out ports
    \-mapi23\ => \-mapi23\,
    \-use.map\ => \-use.map\,
    v0parok => v0parok,
    vm0pari => vm0pari,
    \-vmap0\ => \-vmap0\,
    \-vmap1\ => \-vmap1\,
    \-vmap2\ => \-vmap2\,
    \-vmap3\ => \-vmap3\,
    \-vmap4\ => \-vmap4\,
    vmoparok => vmoparok,
    vpari => vpari
  );
  cadr_vmem1_inst: cadr_vmem1 port map (
      -- in ports
    mapi8 => mapi8,
    mapi9 => mapi9,
    mapi10 => mapi10,
    mapi11 => mapi11,
    mapi12 => mapi12,
    \-vm1wpa\ => \-vm1wpa\,
    \-vma0\ => \-vma0\,
    \-vma1\ => \-vma1\,
    \-vma2\ => \-vma2\,
    \-vma3\ => \-vma3\,
    \-vma4\ => \-vma4\,
    \-vma5\ => \-vma5\,
    \-vma6\ => \-vma6\,
    \-vma7\ => \-vma7\,
    \-vma8\ => \-vma8\,
    \-vma9\ => \-vma9\,
    \-vma10\ => \-vma10\,
    \-vma11\ => \-vma11\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    \-vmap0\ => \-vmap0\,
    \-vmap1\ => \-vmap1\,
    \-vmap2\ => \-vmap2\,
    \-vmap3\ => \-vmap3\,
    \-vmap4\ => \-vmap4\,
      -- out ports
    \-mapi8a\ => \-mapi8a\,
    \-mapi8b\ => \-mapi8b\,
    \-mapi9a\ => \-mapi9a\,
    \-mapi9b\ => \-mapi9b\,
    \-mapi10a\ => \-mapi10a\,
    \-mapi10b\ => \-mapi10b\,
    \-mapi11a\ => \-mapi11a\,
    \-mapi11b\ => \-mapi11b\,
    \-mapi12a\ => \-mapi12a\,
    \-mapi12b\ => \-mapi12b\,
    \-vm1lpar\ => \-vm1lpar\,
    vm1mpar => vm1mpar,
    vm1pari => vm1pari,
    vmap0a => vmap0a,
    vmap1a => vmap1a,
    vmap2a => vmap2a,
    vmap3a => vmap3a,
    vmap4a => vmap4a,
    \-vmo0\ => \-vmo0\,
    \-vmo1\ => \-vmo1\,
    \-vmo2\ => \-vmo2\,
    \-vmo3\ => \-vmo3\,
    \-vmo4\ => \-vmo4\,
    \-vmo5\ => \-vmo5\,
    \-vmo6\ => \-vmo6\,
    \-vmo7\ => \-vmo7\,
    \-vmo8\ => \-vmo8\,
    \-vmo9\ => \-vmo9\,
    \-vmo10\ => \-vmo10\,
    \-vmo11\ => \-vmo11\
  );
  cadr_vmem2_inst: cadr_vmem2 port map (
      -- in ports
    \-mapi8b\ => \-mapi8b\,
    \-mapi9b\ => \-mapi9b\,
    \-mapi10b\ => \-mapi10b\,
    \-mapi11b\ => \-mapi11b\,
    \-mapi12b\ => \-mapi12b\,
    vm1pari => vm1pari,
    \-vm1wpb\ => \-vm1wpb\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    \-vmap0\ => \-vmap0\,
    \-vmap1\ => \-vmap1\,
    \-vmap2\ => \-vmap2\,
    \-vmap3\ => \-vmap3\,
    \-vmap4\ => \-vmap4\,
    \-vmo0\ => \-vmo0\,
    \-vmo1\ => \-vmo1\,
    \-vmo2\ => \-vmo2\,
    \-vmo3\ => \-vmo3\,
    \-vmo4\ => \-vmo4\,
    \-vmo5\ => \-vmo5\,
    \-vmo6\ => \-vmo6\,
    \-vmo7\ => \-vmo7\,
    \-vmo8\ => \-vmo8\,
    \-vmo9\ => \-vmo9\,
    \-vmo10\ => \-vmo10\,
    \-vmo11\ => \-vmo11\,
      -- out ports
    vmap0b => vmap0b,
    vmap1b => vmap1b,
    vmap2b => vmap2b,
    vmap3b => vmap3b,
    vmap4b => vmap4b,
    \-vmo12\ => \-vmo12\,
    \-vmo13\ => \-vmo13\,
    \-vmo14\ => \-vmo14\,
    \-vmo15\ => \-vmo15\,
    \-vmo16\ => \-vmo16\,
    \-vmo17\ => \-vmo17\,
    \-vmo18\ => \-vmo18\,
    \-vmo19\ => \-vmo19\,
    \-vmo20\ => \-vmo20\,
    \-vmo21\ => \-vmo21\,
    \-vmo22\ => \-vmo22\,
    \-vmo23\ => \-vmo23\,
    vmopar => vmopar,
    vmoparck => vmoparck,
    vmoparl => vmoparl,
    vmoparm => vmoparm,
    vmoparodd => vmoparodd
  );
  cadr_vmemdr_inst: cadr_vmemdr port map (
      -- in ports
    hi12 => hi12,
    memstart => memstart,
    \-pfr\ => \-pfr\,
    \-pfw\ => \-pfw\,
    \-srcmap\ => \-srcmap\,
    tse1a => tse1a,
    \-vma0\ => \-vma0\,
    \-vma1\ => \-vma1\,
    \-vma2\ => \-vma2\,
    \-vma3\ => \-vma3\,
    \-vma4\ => \-vma4\,
    \-vma5\ => \-vma5\,
    \-vma6\ => \-vma6\,
    \-vma7\ => \-vma7\,
    \-vmap0\ => \-vmap0\,
    \-vmap1\ => \-vmap1\,
    \-vmap2\ => \-vmap2\,
    \-vmap3\ => \-vmap3\,
    \-vmap4\ => \-vmap4\,
    \-vmo0\ => \-vmo0\,
    \-vmo1\ => \-vmo1\,
    \-vmo2\ => \-vmo2\,
    \-vmo3\ => \-vmo3\,
    \-vmo4\ => \-vmo4\,
    \-vmo5\ => \-vmo5\,
    \-vmo6\ => \-vmo6\,
    \-vmo7\ => \-vmo7\,
    \-vmo8\ => \-vmo8\,
    \-vmo9\ => \-vmo9\,
    \-vmo10\ => \-vmo10\,
    \-vmo11\ => \-vmo11\,
    \-vmo12\ => \-vmo12\,
    \-vmo13\ => \-vmo13\,
    \-vmo14\ => \-vmo14\,
    \-vmo15\ => \-vmo15\,
    \-vmo16\ => \-vmo16\,
    \-vmo17\ => \-vmo17\,
    \-vmo18\ => \-vmo18\,
    \-vmo19\ => \-vmo19\,
    \-vmo20\ => \-vmo20\,
    \-vmo21\ => \-vmo21\,
    \-vmo22\ => \-vmo22\,
    \-vmo23\ => \-vmo23\,
      -- out ports
    \-adrpar\ => \-adrpar\,
    \-lvmo22\ => \-lvmo22\,
    \-lvmo23\ => \-lvmo23\,
    \-mapdrive\ => \-mapdrive\,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    \-pma8\ => \-pma8\,
    \-pma9\ => \-pma9\,
    \-pma10\ => \-pma10\,
    \-pma11\ => \-pma11\,
    \-pma12\ => \-pma12\,
    \-pma13\ => \-pma13\,
    \-pma14\ => \-pma14\,
    \-pma15\ => \-pma15\,
    \-pma16\ => \-pma16\,
    \-pma17\ => \-pma17\,
    \-pma18\ => \-pma18\,
    \-pma19\ => \-pma19\,
    \-pma20\ => \-pma20\,
    \-pma21\ => \-pma21\,
    srcmap => srcmap
  );
  helper_bus_monitor_inst: helper_bus_monitor port map (
      -- in ports
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    aa16 => aa16,
    aa17 => aa17,
    \-aadr0a\ => \-aadr0a\,
    \-aadr1a\ => \-aadr1a\,
    \-aadr2a\ => \-aadr2a\,
    \-aadr3a\ => \-aadr3a\,
    \-aadr4a\ => \-aadr4a\,
    \-aadr5a\ => \-aadr5a\,
    \-aadr6a\ => \-aadr6a\,
    \-aadr7a\ => \-aadr7a\,
    \-aadr8a\ => \-aadr8a\,
    \-aadr9a\ => \-aadr9a\,
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    alu31 => alu31,
    alu32 => alu32,
    aluf0b => aluf0b,
    aluf1b => aluf1b,
    aluf2b => aluf2b,
    aluf3b => aluf3b,
    amem0 => amem0,
    amem1 => amem1,
    amem2 => amem2,
    amem3 => amem3,
    amem4 => amem4,
    amem5 => amem5,
    amem6 => amem6,
    amem7 => amem7,
    amem8 => amem8,
    amem9 => amem9,
    amem10 => amem10,
    amem11 => amem11,
    amem12 => amem12,
    amem13 => amem13,
    amem14 => amem14,
    amem15 => amem15,
    amem16 => amem16,
    amem17 => amem17,
    amem18 => amem18,
    amem19 => amem19,
    amem20 => amem20,
    amem21 => amem21,
    amem22 => amem22,
    amem23 => amem23,
    amem24 => amem24,
    amem25 => amem25,
    amem26 => amem26,
    amem27 => amem27,
    amem28 => amem28,
    amem29 => amem29,
    amem30 => amem30,
    amem31 => amem31,
    dc0 => dc0,
    dc1 => dc1,
    dc2 => dc2,
    dc3 => dc3,
    dc4 => dc4,
    dc5 => dc5,
    dc6 => dc6,
    dc7 => dc7,
    dc8 => dc8,
    dc9 => dc9,
    dpc0 => dpc0,
    dpc1 => dpc1,
    dpc2 => dpc2,
    dpc3 => dpc3,
    dpc4 => dpc4,
    dpc5 => dpc5,
    dpc6 => dpc6,
    dpc7 => dpc7,
    dpc8 => dpc8,
    dpc9 => dpc9,
    dpc10 => dpc10,
    dpc11 => dpc11,
    dpc12 => dpc12,
    dpc13 => dpc13,
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    ipc0 => ipc0,
    ipc1 => ipc1,
    ipc2 => ipc2,
    ipc3 => ipc3,
    ipc4 => ipc4,
    ipc5 => ipc5,
    ipc6 => ipc6,
    ipc7 => ipc7,
    ipc8 => ipc8,
    ipc9 => ipc9,
    ipc10 => ipc10,
    ipc11 => ipc11,
    ipc12 => ipc12,
    ipc13 => ipc13,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir10 => ir10,
    ir11 => ir11,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    ir31 => ir31,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    ir42 => ir42,
    ir43 => ir43,
    ir44 => ir44,
    ir45 => ir45,
    ir46 => ir46,
    ir47 => ir47,
    ir48 => ir48,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lc0 => lc0,
    lc1 => lc1,
    lc2 => lc2,
    lc3 => lc3,
    lc4 => lc4,
    lc5 => lc5,
    lc6 => lc6,
    lc7 => lc7,
    lc8 => lc8,
    lc9 => lc9,
    lc10 => lc10,
    lc11 => lc11,
    lc12 => lc12,
    lc13 => lc13,
    lc14 => lc14,
    lc15 => lc15,
    lc16 => lc16,
    lc17 => lc17,
    lc18 => lc18,
    lc19 => lc19,
    lc20 => lc20,
    lc21 => lc21,
    lc22 => lc22,
    lc23 => lc23,
    lc24 => lc24,
    lc25 => lc25,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    \-madr0a\ => \-madr0a\,
    \-madr1a\ => \-madr1a\,
    \-madr2a\ => \-madr2a\,
    \-madr3a\ => \-madr3a\,
    \-madr4a\ => \-madr4a\,
    mapi8 => mapi8,
    mapi9 => mapi9,
    mapi10 => mapi10,
    mapi11 => mapi11,
    mapi12 => mapi12,
    mapi13 => mapi13,
    mapi14 => mapi14,
    mapi15 => mapi15,
    mapi16 => mapi16,
    mapi17 => mapi17,
    mapi18 => mapi18,
    mapi19 => mapi19,
    mapi20 => mapi20,
    mapi21 => mapi21,
    mapi22 => mapi22,
    mapi23 => mapi23,
    \-md0\ => \-md0\,
    \-md1\ => \-md1\,
    \-md2\ => \-md2\,
    \-md3\ => \-md3\,
    \-md4\ => \-md4\,
    \-md5\ => \-md5\,
    \-md6\ => \-md6\,
    \-md7\ => \-md7\,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-md24\ => \-md24\,
    \-md25\ => \-md25\,
    \-md26\ => \-md26\,
    \-md27\ => \-md27\,
    \-md28\ => \-md28\,
    \-md29\ => \-md29\,
    \-md30\ => \-md30\,
    \-md31\ => \-md31\,
    mem0 => mem0,
    mem1 => mem1,
    mem2 => mem2,
    mem3 => mem3,
    mem4 => mem4,
    mem5 => mem5,
    mem6 => mem6,
    mem7 => mem7,
    mem8 => mem8,
    mem9 => mem9,
    mem10 => mem10,
    mem11 => mem11,
    mem12 => mem12,
    mem13 => mem13,
    mem14 => mem14,
    mem15 => mem15,
    mem16 => mem16,
    mem17 => mem17,
    mem18 => mem18,
    mem19 => mem19,
    mem20 => mem20,
    mem21 => mem21,
    mem22 => mem22,
    mem23 => mem23,
    mem24 => mem24,
    mem25 => mem25,
    mem26 => mem26,
    mem27 => mem27,
    mem28 => mem28,
    mem29 => mem29,
    mem30 => mem30,
    mem31 => mem31,
    mmem0 => mmem0,
    mmem1 => mmem1,
    mmem2 => mmem2,
    mmem3 => mmem3,
    mmem4 => mmem4,
    mmem5 => mmem5,
    mmem6 => mmem6,
    mmem7 => mmem7,
    mmem8 => mmem8,
    mmem9 => mmem9,
    mmem10 => mmem10,
    mmem11 => mmem11,
    mmem12 => mmem12,
    mmem13 => mmem13,
    mmem14 => mmem14,
    mmem15 => mmem15,
    mmem16 => mmem16,
    mmem17 => mmem17,
    mmem18 => mmem18,
    mmem19 => mmem19,
    mmem20 => mmem20,
    mmem21 => mmem21,
    mmem22 => mmem22,
    mmem23 => mmem23,
    mmem24 => mmem24,
    mmem25 => mmem25,
    mmem26 => mmem26,
    mmem27 => mmem27,
    mmem28 => mmem28,
    mmem29 => mmem29,
    mmem30 => mmem30,
    mmem31 => mmem31,
    msk0 => msk0,
    msk1 => msk1,
    msk2 => msk2,
    msk3 => msk3,
    msk4 => msk4,
    msk5 => msk5,
    msk6 => msk6,
    msk7 => msk7,
    msk8 => msk8,
    msk9 => msk9,
    msk10 => msk10,
    msk11 => msk11,
    msk12 => msk12,
    msk13 => msk13,
    msk14 => msk14,
    msk15 => msk15,
    msk16 => msk16,
    msk17 => msk17,
    msk18 => msk18,
    msk19 => msk19,
    msk20 => msk20,
    msk21 => msk21,
    msk22 => msk22,
    msk23 => msk23,
    msk24 => msk24,
    msk25 => msk25,
    msk26 => msk26,
    msk27 => msk27,
    msk28 => msk28,
    msk29 => msk29,
    msk30 => msk30,
    msk31 => msk31,
    npc0 => npc0,
    npc1 => npc1,
    npc2 => npc2,
    npc3 => npc3,
    npc4 => npc4,
    npc5 => npc5,
    npc6 => npc6,
    npc7 => npc7,
    npc8 => npc8,
    npc9 => npc9,
    npc10 => npc10,
    npc11 => npc11,
    npc12 => npc12,
    npc13 => npc13,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    opc0 => opc0,
    opc1 => opc1,
    opc2 => opc2,
    opc3 => opc3,
    opc4 => opc4,
    opc5 => opc5,
    opc6 => opc6,
    opc7 => opc7,
    opc8 => opc8,
    opc9 => opc9,
    opc10 => opc10,
    opc11 => opc11,
    opc12 => opc12,
    opc13 => opc13,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    q0 => q0,
    q1 => q1,
    q2 => q2,
    q3 => q3,
    q4 => q4,
    q5 => q5,
    q6 => q6,
    q7 => q7,
    q8 => q8,
    q9 => q9,
    q10 => q10,
    q11 => q11,
    q12 => q12,
    q13 => q13,
    q14 => q14,
    q15 => q15,
    q16 => q16,
    q17 => q17,
    q18 => q18,
    q19 => q19,
    q20 => q20,
    q21 => q21,
    q22 => q22,
    q23 => q23,
    q24 => q24,
    q25 => q25,
    q26 => q26,
    q27 => q27,
    q28 => q28,
    q29 => q29,
    q30 => q30,
    q31 => q31,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    r7 => r7,
    r8 => r8,
    r9 => r9,
    r10 => r10,
    r11 => r11,
    r12 => r12,
    r13 => r13,
    r14 => r14,
    r15 => r15,
    r16 => r16,
    r17 => r17,
    r18 => r18,
    r19 => r19,
    r20 => r20,
    r21 => r21,
    r22 => r22,
    r23 => r23,
    r24 => r24,
    r25 => r25,
    r26 => r26,
    r27 => r27,
    r28 => r28,
    r29 => r29,
    r30 => r30,
    r31 => r31,
    spc0 => spc0,
    spc1 => spc1,
    spc2 => spc2,
    spc3 => spc3,
    spc4 => spc4,
    spc5 => spc5,
    spc6 => spc6,
    spc7 => spc7,
    spc8 => spc8,
    spc9 => spc9,
    spc10 => spc10,
    spc11 => spc11,
    spc12 => spc12,
    spc13 => spc13,
    spc14 => spc14,
    spc15 => spc15,
    spc16 => spc16,
    spc17 => spc17,
    spc18 => spc18,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15,
    \-vma0\ => \-vma0\,
    \-vma1\ => \-vma1\,
    \-vma2\ => \-vma2\,
    \-vma3\ => \-vma3\,
    \-vma4\ => \-vma4\,
    \-vma5\ => \-vma5\,
    \-vma6\ => \-vma6\,
    \-vma7\ => \-vma7\,
    \-vma8\ => \-vma8\,
    \-vma9\ => \-vma9\,
    \-vma10\ => \-vma10\,
    \-vma11\ => \-vma11\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    \-vma24\ => \-vma24\,
    \-vma25\ => \-vma25\,
    \-vma26\ => \-vma26\,
    \-vma27\ => \-vma27\,
    \-vma28\ => \-vma28\,
    \-vma29\ => \-vma29\,
    \-vma30\ => \-vma30\,
    \-vma31\ => \-vma31\,
    wadr0 => wadr0,
    wadr1 => wadr1,
    wadr2 => wadr2,
    wadr3 => wadr3,
    wadr4 => wadr4,
    wadr5 => wadr5,
    wadr6 => wadr6,
    wadr7 => wadr7,
    wadr8 => wadr8,
    wadr9 => wadr9
  );
  helper_required_signals_inst: helper_required_signals port map (
      -- in ports
    \bus.power.reset l\ => \bus.power.reset l\,
    \-bus.reset\ => \-bus.reset\,
    mclk7 => mclk7,
      -- out ports
    \-boot1\ => \-boot1\,
    \-busint.lm.reset\ => \-busint.lm.reset\,
    \-dbread\ => \-dbread\,
    \-dbwrite\ => \-dbwrite\,
    eadr0 => eadr0,
    eadr1 => eadr1,
    eadr2 => eadr2,
    eadr3 => eadr3,
    \-halt\ => \-halt\,
    \lm drive enb\ => \lm drive enb\
  );
end architecture;
