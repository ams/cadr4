library ieee;
use ieee.std_logic_1164.all;

entity cadr_npc is
  port (
    ipc13   : out std_logic;
    pc13    : out std_logic;
    ipc12   : out std_logic;
    pc12    : out std_logic;
    pccry11 : out std_logic;
    ipc9    : out std_logic;
    pc9     : out std_logic;
    ipc8    : out std_logic;
    pc8     : out std_logic;
    pccry7  : out std_logic;
    ipc11   : out std_logic;
    pc11    : out std_logic;
    ipc10   : out std_logic;
    pc10    : out std_logic;
    ipc5    : out std_logic;
    pc5     : out std_logic;
    pc4     : out std_logic;
    pccry3  : out std_logic;
    ipc7    : out std_logic;
    pc7     : out std_logic;
    ipc6    : out std_logic;
    pc6     : out std_logic;
    ipc1    : out std_logic;
    pc1     : out std_logic;
    ipc0    : out std_logic;
    pc0     : out std_logic;
    ipc3    : out std_logic;
    pc3     : out std_logic;
    ipc2    : out std_logic;
    pc2     : out std_logic;
    trapb   : in  std_logic;
    pcs1    : in  std_logic;
    dpc3    : out std_logic;
    ir15    : in  std_logic;
    spc3    : out std_logic;
    npc3    : out std_logic;
    npc2    : out std_logic;
    spc2    : out std_logic;
    ir14    : in  std_logic;
    dpc2    : out std_logic;
    pcs0    : in  std_logic;
    dpc1    : out std_logic;
    ir13    : in  std_logic;
    spc1a   : in  std_logic;
    npc1    : out std_logic;
    npc0    : out std_logic;
    spc0    : out std_logic;
    ir12    : in  std_logic;
    dpc0    : out std_logic;
    npc13   : out std_logic;
    npc12   : out std_logic;
    clk4b   : in  std_logic;
    npc11   : out std_logic;
    npc10   : out std_logic;
    npc9    : out std_logic;
    npc8    : out std_logic;
    npc7    : out std_logic;
    npc6    : out std_logic;
    npc5    : out std_logic;
    npc4    : out std_logic;
    trapa   : in  std_logic;
    dpc13   : out std_logic;
    ir25    : in  std_logic;
    spc13   : out std_logic;
    spc12   : out std_logic;
    ir24    : in  std_logic;
    dpc12   : out std_logic;
    dpc11   : out std_logic;
    ir23    : in  std_logic;
    spc11   : out std_logic;
    spc10   : out std_logic;
    ir22    : in  std_logic;
    dpc10   : out std_logic;
    dpc9    : out std_logic;
    ir21    : in  std_logic;
    spc9    : out std_logic;
    spc8    : out std_logic;
    ir20    : in  std_logic;
    dpc8    : out std_logic;
    dpc7    : out std_logic;
    ir19    : in  std_logic;
    spc7    : out std_logic;
    spc6    : out std_logic;
    ir18    : in  std_logic;
    dpc6    : out std_logic;
    dpc5    : out std_logic;
    ir17    : in  std_logic;
    spc5    : out std_logic;
    spc4    : out std_logic;
    ir16    : in  std_logic;
    dpc4    : in  std_logic;
    ipc4    : out std_logic
    );
end;
