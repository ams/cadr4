library ieee;
use ieee.std_logic_1164.all;

entity cadr_opcd is
  port (
    \-srcdc\        : in     std_logic;
    \-srcopc\       : in     std_logic;
    \-srcpdlidx\    : in     std_logic;
    \-srcpdlptr\    : in     std_logic;
    dc0             : in     std_logic;
    dc1             : in     std_logic;
    dc2             : in     std_logic;
    dc3             : in     std_logic;
    dc4             : in     std_logic;
    dc5             : in     std_logic;
    dc6             : in     std_logic;
    dc7             : in     std_logic;
    dc8             : in     std_logic;
    dc9             : in     std_logic;
    opc0            : in     std_logic;
    opc1            : in     std_logic;
    opc10           : in     std_logic;
    opc11           : in     std_logic;
    opc12           : in     std_logic;
    opc13           : in     std_logic;
    opc2            : in     std_logic;
    opc3            : in     std_logic;
    opc4            : in     std_logic;
    opc5            : in     std_logic;
    opc6            : in     std_logic;
    opc7            : in     std_logic;
    opc8            : in     std_logic;
    opc9            : in     std_logic;
    tse1b           : in     std_logic;
    \-opcdrive\     : out    std_logic;
    \-zero16.drive\ : out    std_logic;
    \zero12.drive\  : out    std_logic;
    \zero16.drive\  : out    std_logic;
    dcdrive         : out    std_logic;
    mf0             : out    std_logic;
    mf1             : out    std_logic;
    mf10            : out    std_logic;
    mf11            : out    std_logic;
    mf12            : out    std_logic;
    mf13            : out    std_logic;
    mf14            : out    std_logic;
    mf15            : out    std_logic;
    mf16            : out    std_logic;
    mf17            : out    std_logic;
    mf18            : out    std_logic;
    mf19            : out    std_logic;
    mf2             : out    std_logic;
    mf20            : out    std_logic;
    mf21            : out    std_logic;
    mf22            : out    std_logic;
    mf23            : out    std_logic;
    mf24            : out    std_logic;
    mf25            : out    std_logic;
    mf26            : out    std_logic;
    mf27            : out    std_logic;
    mf28            : out    std_logic;
    mf29            : out    std_logic;
    mf3             : out    std_logic;
    mf30            : out    std_logic;
    mf31            : out    std_logic;
    mf4             : out    std_logic;
    mf5             : out    std_logic;
    mf6             : out    std_logic;
    mf7             : out    std_logic;
    mf8             : out    std_logic;
    mf9             : out    std_logic;
    zero16          : out    std_logic
  );
end entity cadr_opcd;
