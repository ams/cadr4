library ieee;
use ieee.std_logic_1164.all;

package utilities is

end package utilities;

package body utilities is

end package body utilities;
