library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn7408_tb is
end sn7408_tb;

architecture testbench of sn7408_tb is

begin

--  uut : sn7408 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
