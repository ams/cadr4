library ieee;
use ieee.std_logic_1164.all;

entity cadr_shift1 is
  port (
    \-s4\           : in     std_logic;
    m13             : in     std_logic;
    m14             : in     std_logic;
    m15             : in     std_logic;
    m16             : in     std_logic;
    m17             : in     std_logic;
    m18             : in     std_logic;
    m19             : in     std_logic;
    m20             : in     std_logic;
    m21             : in     std_logic;
    m22             : in     std_logic;
    m23             : in     std_logic;
    m24             : in     std_logic;
    m25             : in     std_logic;
    m26             : in     std_logic;
    m27             : in     std_logic;
    m28             : in     std_logic;
    m29             : in     std_logic;
    m30             : in     std_logic;
    m31             : in     std_logic;
    s0              : in     std_logic;
    s1              : in     std_logic;
    s2b             : in     std_logic;
    s3b             : in     std_logic;
    s4              : in     std_logic;
    sa0             : in     std_logic;
    sa1             : in     std_logic;
    sa10            : in     std_logic;
    sa11            : in     std_logic;
    sa12            : in     std_logic;
    sa13            : in     std_logic;
    sa14            : in     std_logic;
    sa15            : in     std_logic;
    sa2             : in     std_logic;
    sa3             : in     std_logic;
    sa4             : in     std_logic;
    sa5             : in     std_logic;
    sa6             : in     std_logic;
    sa7             : in     std_logic;
    sa8             : in     std_logic;
    sa9             : in     std_logic;
    r16             : out    std_logic;
    r17             : out    std_logic;
    r18             : out    std_logic;
    r19             : out    std_logic;
    r20             : out    std_logic;
    r21             : out    std_logic;
    r22             : out    std_logic;
    r23             : out    std_logic;
    r24             : out    std_logic;
    r25             : out    std_logic;
    r26             : out    std_logic;
    r27             : out    std_logic;
    r28             : out    std_logic;
    r29             : out    std_logic;
    r30             : out    std_logic;
    r31             : out    std_logic;
    sa16            : out    std_logic;
    sa17            : out    std_logic;
    sa18            : out    std_logic;
    sa19            : out    std_logic;
    sa20            : out    std_logic;
    sa21            : out    std_logic;
    sa22            : out    std_logic;
    sa23            : out    std_logic;
    sa24            : out    std_logic;
    sa25            : out    std_logic;
    sa26            : out    std_logic;
    sa27            : out    std_logic;
    sa28            : out    std_logic;
    sa29            : out    std_logic;
    sa30            : out    std_logic;
    sa31            : out    std_logic
  );
end entity;
