-- 4096 X 1 Bt Static RAM
-- Intel 2147H
-- doc/ttl/d2147.pdf

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity d2147 is
  port (
    a0   : in  std_logic := 'H';
    a1   : in  std_logic := 'H';
    a2   : in  std_logic := 'H';
    a3   : in  std_logic := 'H';
    a4   : in  std_logic := 'H';
    a5   : in  std_logic := 'H';
    a6   : in  std_logic := 'H';
    a7   : in  std_logic := 'H';
    a8   : in  std_logic := 'H';
    a9   : in  std_logic := 'H';
    a10  : in  std_logic := 'H';
    a11  : in  std_logic := 'H';
    ce_n : in  std_logic := 'H';
    di   : in  std_logic := 'H';
    we_n : in  std_logic := 'H';
    do   : out std_logic
    );
end entity;

architecture ttl of d2147 is
  type ram_t is array (0 to 4095) of std_logic;
  signal ram : ram_t := (others => '0');
begin
  process (all)
    variable addr : unsigned(11 downto 0);
  begin
    if to_x01(ce_n) = '0' then
      addr := (a11, a10, a9, a8, a7, a6, a5, a4, a3, a2, a1, a0);
      if is_x(addr) then
        if to_x01(we_n) = '1' then
          do <= 'X';
        end if;
      else
        if to_x01(we_n) = '0' then
          ram(to_integer(addr)) <= di;
        elsif to_x01(we_n) = '1' then
          do <= ram(to_integer(addr));
        else
          -- do nothing
        end if;
      end if;
    elsif to_x01(ce_n) = '1' then
      do <= 'Z';
    else
      do <= 'X';
    end if;
  end process;
end architecture;
