-- CADR1_BUSSEL
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_bussel is
  port (
    \-ub16_bus\ : in std_logic;
    \-ub32_bus\ : in std_logic;
    bus0 : out std_logic;
    bus1 : out std_logic;
    bus10 : out std_logic;
    bus11 : out std_logic;
    bus12 : out std_logic;
    bus13 : out std_logic;
    bus14 : out std_logic;
    bus15 : out std_logic;
    bus16 : out std_logic;
    bus17 : out std_logic;
    bus18 : out std_logic;
    bus19 : out std_logic;
    bus2 : out std_logic;
    bus20 : out std_logic;
    bus21 : out std_logic;
    bus22 : out std_logic;
    bus23 : out std_logic;
    bus24 : out std_logic;
    bus25 : out std_logic;
    bus26 : out std_logic;
    bus27 : out std_logic;
    bus28 : out std_logic;
    bus29 : out std_logic;
    bus3 : out std_logic;
    bus30 : out std_logic;
    bus31 : out std_logic;
    bus4 : out std_logic;
    bus5 : out std_logic;
    bus6 : out std_logic;
    bus7 : out std_logic;
    bus8 : out std_logic;
    bus9 : out std_logic;
    udi0 : in std_logic;
    udi1 : in std_logic;
    udi10 : in std_logic;
    udi11 : in std_logic;
    udi12 : in std_logic;
    udi13 : in std_logic;
    udi14 : in std_logic;
    udi15 : in std_logic;
    udi2 : in std_logic;
    udi3 : in std_logic;
    udi4 : in std_logic;
    udi5 : in std_logic;
    udi6 : in std_logic;
    udi7 : in std_logic;
    udi8 : in std_logic;
    udi9 : in std_logic;
    wbuf0 : in std_logic;
    wbuf1 : in std_logic;
    wbuf10 : in std_logic;
    wbuf11 : in std_logic;
    wbuf12 : in std_logic;
    wbuf13 : in std_logic;
    wbuf14 : in std_logic;
    wbuf15 : in std_logic;
    wbuf2 : in std_logic;
    wbuf3 : in std_logic;
    wbuf4 : in std_logic;
    wbuf5 : in std_logic;
    wbuf6 : in std_logic;
    wbuf7 : in std_logic;
    wbuf8 : in std_logic;
    wbuf9 : in std_logic
  );
end entity;
