library ieee;
use ieee.std_logic_1164.all;

entity cadr_spy1 is
  port (
    \-spy.obl\ : out std_logic;
    ob7        : in  std_logic;
    spy0       : out std_logic;
    ob6        : in  std_logic;
    spy1       : out std_logic;
    ob5        : in  std_logic;
    spy2       : out std_logic;
    ob4        : in  std_logic;
    spy3       : out std_logic;
    ob3        : in  std_logic;
    spy4       : out std_logic;
    ob2        : in  std_logic;
    spy5       : out std_logic;
    ob1        : in  std_logic;
    spy6       : out std_logic;
    ob0        : in  std_logic;
    spy7       : out std_logic;
    ob15       : in  std_logic;
    spy8       : out std_logic;
    ob14       : in  std_logic;
    spy9       : out std_logic;
    ob13       : in  std_logic;
    spy10      : out std_logic;
    ob12       : in  std_logic;
    spy11      : out std_logic;
    ob11       : in  std_logic;
    spy12      : out std_logic;
    ob10       : in  std_logic;
    spy13      : out std_logic;
    ob9        : in  std_logic;
    spy14      : out std_logic;
    ob8        : in  std_logic;
    spy15      : out std_logic;
    \-spy.obh\ : in  std_logic;
    ob23       : in  std_logic;
    ob22       : in  std_logic;
    ob21       : in  std_logic;
    ob20       : in  std_logic;
    ob19       : in  std_logic;
    ob18       : in  std_logic;
    ob17       : in  std_logic;
    ob16       : in  std_logic;
    ob31       : in  std_logic;
    ob30       : in  std_logic;
    ob29       : in  std_logic;
    ob28       : in  std_logic;
    ob27       : in  std_logic;
    ob26       : in  std_logic;
    ob25       : in  std_logic;
    ob24       : in  std_logic;
    \-spy.irl\ : in  std_logic;
    ir7        : in  std_logic;
    ir6        : in  std_logic;
    ir5        : in  std_logic;
    ir4        : in  std_logic;
    ir3        : in  std_logic;
    ir2        : in  std_logic;
    ir1        : in  std_logic;
    ir0        : in  std_logic;
    ir15       : in  std_logic;
    ir14       : in  std_logic;
    ir13       : in  std_logic;
    ir12       : in  std_logic;
    ir11       : in  std_logic;
    ir10       : in  std_logic;
    ir9        : in  std_logic;
    ir8        : in  std_logic;
    \-spy.irh\ : in  std_logic;
    ir47       : in  std_logic;
    ir46       : in  std_logic;
    ir45       : in  std_logic;
    ir44       : in  std_logic;
    ir43       : in  std_logic;
    ir42       : in  std_logic;
    ir41       : in  std_logic;
    ir40       : in  std_logic;
    ir39       : in  std_logic;
    ir38       : in  std_logic;
    ir37       : in  std_logic;
    ir36       : in  std_logic;
    ir35       : in  std_logic;
    ir34       : in  std_logic;
    ir33       : in  std_logic;
    ir32       : in  std_logic;
    \-spy.irm\ : in  std_logic;
    ir31       : in  std_logic;
    ir30       : in  std_logic;
    ir29       : in  std_logic;
    ir28       : in  std_logic;
    ir27       : in  std_logic;
    ir26       : in  std_logic;
    ir25       : in  std_logic;
    ir24       : in  std_logic;
    ir23       : in  std_logic;
    ir22       : in  std_logic;
    ir21       : in  std_logic;
    ir20       : in  std_logic;
    ir19       : in  std_logic;
    ir18       : in  std_logic;
    ir17       : in  std_logic;
    ir16       : in  std_logic
    );
end;
