-- PDL1 -- PDL BUFFER RIGHT

library work;
use work.dip.all;
use work.misc.all;

architecture behv of cadr_pdl1 is
begin
pdl1_4c21 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl13, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpb\, p15 => l13);
pdl1_4c23 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl12, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpb\, p15 => l12);
pdl1_4c24 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl11, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpb\, p15 => l11);
pdl1_4c25 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl10, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l10);
pdl1_4c26 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl4, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l4);
pdl1_4c27 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl3, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l3);
pdl1_4c28 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl2, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l2);
pdl1_4c29 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl1, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l1);
pdl1_4c30 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl0, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l0);
pdl1_4d23 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl15, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpb\, p15 => l15);
pdl1_4d25 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl14, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpb\, p15 => l14);
pdl1_4d26 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl9, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l9);
pdl1_4d27 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl8, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l8);
pdl1_4d28 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl7, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l7);
pdl1_4d29 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl6, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l6);
pdl1_4d30 : dip_93425a port map (p1 => gnd, p2 => \-pdla0a\, p3 => \-pdla1a\, p4 => \-pdla2a\, p5 => \-pdla3a\, p6 => \-pdla4a\, p7 => pdl5, p9 => \-pdla5a\, p10 => \-pdla6a\, p11 => \-pdla7a\, p12 => \-pdla8a\, p13 => \-pdla9a\, p14 => \-pwpc\, p15 => l5);
end architecture;
