library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_shift1 is
  port (
    m21   : in  std_logic;
    m22   : in  std_logic;
    m23   : in  std_logic;
    m24   : in  std_logic;
    m25   : in  std_logic;
    m26   : in  std_logic;
    m27   : in  std_logic;
    s1    : in  std_logic;
    s0    : in  std_logic;
    sa27  : out std_logic;
    sa26  : out std_logic;
    gnd   : in  std_logic;
    sa25  : out std_logic;
    sa24  : out std_logic;
    m13   : in  std_logic;
    m14   : in  std_logic;
    m15   : in  std_logic;
    m16   : in  std_logic;
    m17   : in  std_logic;
    m18   : in  std_logic;
    m19   : in  std_logic;
    sa19  : out std_logic;
    sa18  : out std_logic;
    sa17  : out std_logic;
    sa16  : out std_logic;
    m28   : in  std_logic;
    m29   : in  std_logic;
    m30   : in  std_logic;
    m31   : in  std_logic;
    sa31  : out std_logic;
    sa30  : out std_logic;
    sa29  : out std_logic;
    sa28  : out std_logic;
    m20   : in  std_logic;
    sa23  : out std_logic;
    sa22  : out std_logic;
    sa21  : out std_logic;
    sa20  : out std_logic;
    sa2   : in  std_logic;
    sa6   : in  std_logic;
    sa10  : in  std_logic;
    sa14  : in  std_logic;
    s3b   : in  std_logic;
    s2b   : in  std_logic;
    r30   : out std_logic;
    r26   : out std_logic;
    \-s4\ : in  std_logic;
    r22   : out std_logic;
    r18   : out std_logic;
    s4    : in  std_logic;
    sa3   : in  std_logic;
    sa7   : in  std_logic;
    sa11  : in  std_logic;
    sa15  : in  std_logic;
    r31   : out std_logic;
    r27   : out std_logic;
    r23   : out std_logic;
    r19   : out std_logic;
    sa0   : in  std_logic;
    sa4   : in  std_logic;
    sa8   : in  std_logic;
    sa12  : in  std_logic;
    r28   : out std_logic;
    r24   : out std_logic;
    r20   : out std_logic;
    r16   : out std_logic;
    sa1   : in  std_logic;
    sa5   : in  std_logic;
    sa9   : in  std_logic;
    sa13  : in  std_logic;
    r29   : out std_logic;
    r25   : out std_logic;
    r21   : out std_logic;
    r17   : out std_logic);
end;

architecture ttl of cadr_shift1 is
begin
  shift1_2c01 : am25s10 port map(i_3 => m21, i_2 => m22, i_1 => m23, i0 => m24, i1 => m25, i2 => m26, i3 => m27, sel1 => s1, sel0 => s0, o3 => sa27, o2 => sa26, ce_n => gnd, o1 => sa25, o0 => sa24);
  shift1_2c06 : am25s10 port map(i_3 => m13, i_2 => m14, i_1 => m15, i0 => m16, i1 => m17, i2 => m18, i3 => m19, sel1 => s1, sel0 => s0, o3 => sa19, o2 => sa18, ce_n => gnd, o1 => sa17, o0 => sa16);
  shift1_2d05 : am25s10 port map(i_3 => m25, i_2 => m26, i_1 => m27, i0 => m28, i1 => m29, i2 => m30, i3 => m31, sel1 => s1, sel0 => s0, o3 => sa31, o2 => sa30, ce_n => gnd, o1 => sa29, o0 => sa28);
  shift1_2d10 : am25s10 port map(i_3 => m17, i_2 => m18, i_1 => m19, i0 => m20, i1 => m21, i2 => m22, i3 => m23, sel1 => s1, sel0 => s0, o3 => sa23, o2 => sa22, ce_n => gnd, o1 => sa21, o0 => sa20);
  shift1_2e01 : am25s10 port map(i_3 => sa22, i_2 => sa26, i_1 => sa30, i0 => sa2, i1 => sa6, i2 => sa10, i3 => sa14, sel1 => s3b, sel0 => s2b, o3 => r30, o2 => r26, ce_n => \-s4\, o1 => r22, o0 => r18);
  shift1_2e02 : am25s10 port map(i_3 => sa6, i_2 => sa10, i_1 => sa14, i0 => sa18, i1 => sa22, i2 => sa26, i3 => sa30, sel1 => s3b, sel0 => s2b, o3 => r30, o2 => r26, ce_n => s4, o1 => r22, o0 => r18);
  shift1_2e03 : am25s10 port map(i_3 => sa23, i_2 => sa27, i_1 => sa31, i0 => sa3, i1 => sa7, i2 => sa11, i3 => sa15, sel1 => s3b, sel0 => s2b, o3 => r31, o2 => r27, ce_n => \-s4\, o1 => r23, o0 => r19);
  shift1_2e04 : am25s10 port map(i_3 => sa7, i_2 => sa11, i_1 => sa15, i0 => sa19, i1 => sa23, i2 => sa27, i3 => sa31, sel1 => s3b, sel0 => s2b, o3 => r31, o2 => r27, ce_n => s4, o1 => r23, o0 => r19);
  shift1_2e06 : am25s10 port map(i_3 => sa20, i_2 => sa24, i_1 => sa28, i0 => sa0, i1 => sa4, i2 => sa8, i3 => sa12, sel1 => s3b, sel0 => s2b, o3 => r28, o2 => r24, ce_n => \-s4\, o1 => r20, o0 => r16);
  shift1_2e07 : am25s10 port map(i_3 => sa4, i_2 => sa8, i_1 => sa12, i0 => sa16, i1 => sa20, i2 => sa24, i3 => sa28, sel1 => s3b, sel0 => s2b, o3 => r28, o2 => r24, ce_n => s4, o1 => r20, o0 => r16);
  shift1_2e08 : am25s10 port map(i_3 => sa21, i_2 => sa25, i_1 => sa29, i0 => sa1, i1 => sa5, i2 => sa9, i3 => sa13, sel1 => s3b, sel0 => s2b, o3 => r29, o2 => r25, ce_n => \-s4\, o1 => r21, o0 => r17);
  shift1_2e09 : am25s10 port map(i_3 => sa5, i_2 => sa9, i_1 => sa13, i0 => sa17, i1 => sa21, i2 => sa25, i3 => sa29, sel1 => s3b, sel0 => s2b, o3 => r29, o2 => r25, ce_n => s4, o1 => r21, o0 => r17);
end architecture;
