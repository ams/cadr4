library ieee;
use ieee.std_logic_1164.all;

entity cadr1_uprior is
  port (
    \-clk\          : in     std_logic;
    \-disable int grant\ : in     std_logic;
    \-local enable\ : in     std_logic;
    \-npg in\       : in     std_logic;
    \-npg out\      : in     std_logic;
    \-ub br4\       : in     std_logic;
    \-ub br5\       : in     std_logic;
    \-ub br6\       : in     std_logic;
    \-ub br7\       : in     std_logic;
    \-ub init\      : in     std_logic;
    \-ub intr\      : in     std_logic;
    \-ub npr\       : in     std_logic;
    \bus req\       : in     std_logic;
    \grant timeout\ : in     std_logic;
    \hi 1-14\       : in     std_logic;
    \local enable\  : in     std_logic;
    \sack in\       : in     std_logic;
    \unibus init in\ : in     std_logic;
    \unibus intr in\ : in     std_logic;
    br4             : in     std_logic;
    br5             : in     std_logic;
    br6             : in     std_logic;
    br7             : in     std_logic;
    level0          : in     std_logic;
    level1          : in     std_logic;
    npr             : in     std_logic;
    reset           : in     std_logic;
    \-bg4o\         : inout  std_logic;
    \-bg5o\         : inout  std_logic;
    \-bg6o\         : inout  std_logic;
    \-bg7o\         : inout  std_logic;
    \-clear grant\  : inout  std_logic;
    \-npgo\         : inout  std_logic;
    \any grant dlyd\ : inout  std_logic;
    \any grant\     : inout  std_logic;
    \ub npg in\     : inout  std_logic;
    \ub npg out\    : inout  std_logic;
    bg4p            : inout  std_logic;
    bg5p            : inout  std_logic;
    bg6p            : inout  std_logic;
    bg7p            : inout  std_logic;
    br4d            : inout  std_logic;
    br5d            : inout  std_logic;
    br6d            : inout  std_logic;
    br7d            : inout  std_logic;
    npgp            : inout  std_logic;
    nprd            : inout  std_logic;
    sackd           : inout  std_logic;
    \-any grant dlyd\ : out    std_logic;
    \any int grant\ : out    std_logic;
    \ub bg4 in\     : out    std_logic;
    \ub bg5 in\     : out    std_logic;
    \ub bg6 in\     : out    std_logic;
    \ub bg7 in\     : out    std_logic;
    bg4o            : out    std_logic;
    bg5o            : out    std_logic;
    bg6o            : out    std_logic;
    bg7o            : out    std_logic;
    npgo            : out    std_logic
  );
end entity cadr1_uprior;
