library ieee;
use ieee.std_logic_1164.all;

entity cadr_ipar is
  port (
    imodd           : in     std_logic;
    ir0             : in     std_logic;
    ir1             : in     std_logic;
    ir10            : in     std_logic;
    ir11            : in     std_logic;
    ir12            : in     std_logic;
    ir13            : in     std_logic;
    ir14            : in     std_logic;
    ir15            : in     std_logic;
    ir16            : in     std_logic;
    ir17            : in     std_logic;
    ir18            : in     std_logic;
    ir19            : in     std_logic;
    ir2             : in     std_logic;
    ir20            : in     std_logic;
    ir21            : in     std_logic;
    ir22            : in     std_logic;
    ir23            : in     std_logic;
    ir24            : in     std_logic;
    ir25            : in     std_logic;
    ir26            : in     std_logic;
    ir27            : in     std_logic;
    ir28            : in     std_logic;
    ir29            : in     std_logic;
    ir3             : in     std_logic;
    ir30            : in     std_logic;
    ir31            : in     std_logic;
    ir32            : in     std_logic;
    ir33            : in     std_logic;
    ir34            : in     std_logic;
    ir35            : in     std_logic;
    ir36            : in     std_logic;
    ir37            : in     std_logic;
    ir38            : in     std_logic;
    ir39            : in     std_logic;
    ir4             : in     std_logic;
    ir40            : in     std_logic;
    ir41            : in     std_logic;
    ir42            : in     std_logic;
    ir43            : in     std_logic;
    ir44            : in     std_logic;
    ir45            : in     std_logic;
    ir46            : in     std_logic;
    ir47            : in     std_logic;
    ir48            : in     std_logic;
    ir5             : in     std_logic;
    ir6             : in     std_logic;
    ir7             : in     std_logic;
    ir8             : in     std_logic;
    ir9             : in     std_logic;
    ipar0           : out    std_logic;
    ipar1           : out    std_logic;
    ipar2           : out    std_logic;
    ipar3           : out    std_logic;
    iparity         : out    std_logic;
    iparok          : out    std_logic
  );
end entity cadr_ipar;
