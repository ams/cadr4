library ieee;
use ieee.std_logic_1164.all;

entity cadr_lc is
  port (
    \-lcdrive\          : out std_logic;
    needfetch           : in  std_logic;
    mf24                : out std_logic;
    gnd                 : in  std_logic;
    mf25                : out std_logic;
    \lc byte mode\      : in  std_logic;
    mf26                : out std_logic;
    \prog.unibus.reset\ : in  std_logic;
    mf27                : out std_logic;
    \int.enable\        : in  std_logic;
    mf28                : out std_logic;
    \sequence.break\    : in  std_logic;
    mf29                : out std_logic;
    lc25                : out std_logic;
    mf30                : out std_logic;
    lc24                : out std_logic;
    mf31                : out std_logic;
    lcdrive             : out std_logic;
    srclc               : out std_logic;
    tse1a               : in  std_logic;
    lc7                 : out std_logic;
    mf0                 : out std_logic;
    lc6                 : out std_logic;
    mf1                 : out std_logic;
    lc5                 : out std_logic;
    mf2                 : out std_logic;
    lc4                 : out std_logic;
    mf3                 : out std_logic;
    lc3                 : in  std_logic;
    mf4                 : out std_logic;
    lc2                 : in  std_logic;
    mf5                 : out std_logic;
    lc1                 : in  std_logic;
    mf6                 : out std_logic;
    lc0b                : in  std_logic;
    mf7                 : out std_logic;
    lc23                : out std_logic;
    mf16                : out std_logic;
    lc22                : out std_logic;
    mf17                : out std_logic;
    lc21                : out std_logic;
    mf18                : out std_logic;
    lc20                : out std_logic;
    mf19                : out std_logic;
    lc19                : out std_logic;
    mf20                : out std_logic;
    lc18                : out std_logic;
    mf21                : out std_logic;
    lc17                : out std_logic;
    mf22                : out std_logic;
    lc16                : out std_logic;
    mf23                : out std_logic;
    lc15                : out std_logic;
    mf8                 : out std_logic;
    lc14                : out std_logic;
    mf9                 : out std_logic;
    lc13                : out std_logic;
    mf10                : out std_logic;
    lc12                : out std_logic;
    mf11                : out std_logic;
    lc11                : out std_logic;
    mf12                : out std_logic;
    lc10                : out std_logic;
    mf13                : out std_logic;
    lc9                 : out std_logic;
    mf14                : out std_logic;
    lc8                 : out std_logic;
    mf15                : out std_logic;
    hi11                : in  std_logic;
    clk1a               : in  std_logic;
    ob20                : in  std_logic;
    ob21                : in  std_logic;
    ob22                : in  std_logic;
    ob23                : in  std_logic;
    \-destlc\           : in  std_logic;
    \-lcry19\           : out std_logic;
    \-lcry23\           : out std_logic;
    ob16                : in  std_logic;
    ob17                : in  std_logic;
    ob18                : in  std_logic;
    ob19                : in  std_logic;
    \-lcry15\           : out std_logic;
    clk2a               : in  std_logic;
    ob12                : in  std_logic;
    ob13                : in  std_logic;
    ob14                : in  std_logic;
    ob15                : in  std_logic;
    \-lcry11\           : out std_logic;
    clk2c               : in  std_logic;
    ob8                 : in  std_logic;
    ob9                 : in  std_logic;
    ob10                : in  std_logic;
    ob11                : in  std_logic;
    \-srclc\            : in  std_logic;
    ob24                : in  std_logic;
    ob25                : in  std_logic;
    ob4                 : in  std_logic;
    ob5                 : in  std_logic;
    ob6                 : in  std_logic;
    ob7                 : in  std_logic;
    \-lcry3\            : in  std_logic;
    \-lcry7\            : out std_logic
    );
end;
