library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;

entity sn7432_tb is
end sn7432_tb;

architecture testbench of sn7432_tb is

begin

--  uut : sn7432 port map(
--    );

  process
  begin
    wait for 5 ns;

    wait;
  end process;

end testbench;
