library ieee;
use ieee.std_logic_1164.all;

entity cadr1_xd is
  port (
    \-xbus ignpar\  : in     std_logic;
    \-xbus par\     : in     std_logic;
    \-xbus wr\      : in     std_logic;
    \-xbus0\        : in     std_logic;
    \-xbus10\       : in     std_logic;
    \-xbus11\       : in     std_logic;
    \-xbus12\       : in     std_logic;
    \-xbus13\       : in     std_logic;
    \-xbus14\       : in     std_logic;
    \-xbus15\       : in     std_logic;
    \-xbus16\       : in     std_logic;
    \-xbus17\       : in     std_logic;
    \-xbus18\       : in     std_logic;
    \-xbus19\       : in     std_logic;
    \-xbus1\        : in     std_logic;
    \-xbus20\       : in     std_logic;
    \-xbus21\       : in     std_logic;
    \-xbus22\       : in     std_logic;
    \-xbus23\       : in     std_logic;
    \-xbus24\       : in     std_logic;
    \-xbus25\       : in     std_logic;
    \-xbus26\       : in     std_logic;
    \-xbus27\       : in     std_logic;
    \-xbus28\       : in     std_logic;
    \-xbus29\       : in     std_logic;
    \-xbus2\        : in     std_logic;
    \-xbus30\       : in     std_logic;
    \-xbus31\       : in     std_logic;
    \-xbus3\        : in     std_logic;
    \-xbus4\        : in     std_logic;
    \-xbus5\        : in     std_logic;
    \-xbus6\        : in     std_logic;
    \-xbus7\        : in     std_logic;
    \-xbus8\        : in     std_logic;
    \-xbus9\        : in     std_logic;
    \-xdrive\       : in     std_logic;
    \hi 15-30\      : in     std_logic;
    \xbus ignpar in\ : in     std_logic;
    \xbus par in\   : in     std_logic;
    \xbus par out\  : in     std_logic;
    bus0            : in     std_logic;
    bus1            : in     std_logic;
    bus10           : in     std_logic;
    bus11           : in     std_logic;
    bus12           : in     std_logic;
    bus13           : in     std_logic;
    bus14           : in     std_logic;
    bus15           : in     std_logic;
    bus16           : in     std_logic;
    bus17           : in     std_logic;
    bus18           : in     std_logic;
    bus19           : in     std_logic;
    bus2            : in     std_logic;
    bus20           : in     std_logic;
    bus21           : in     std_logic;
    bus22           : in     std_logic;
    bus23           : in     std_logic;
    bus24           : in     std_logic;
    bus25           : in     std_logic;
    bus26           : in     std_logic;
    bus27           : in     std_logic;
    bus28           : in     std_logic;
    bus29           : in     std_logic;
    bus3            : in     std_logic;
    bus30           : in     std_logic;
    bus31           : in     std_logic;
    bus4            : in     std_logic;
    bus5            : in     std_logic;
    bus6            : in     std_logic;
    bus7            : in     std_logic;
    bus8            : in     std_logic;
    bus9            : in     std_logic;
    xdi0            : in     std_logic;
    xdi1            : in     std_logic;
    xdi10           : in     std_logic;
    xdi11           : in     std_logic;
    xdi12           : in     std_logic;
    xdi13           : in     std_logic;
    xdi14           : in     std_logic;
    xdi15           : in     std_logic;
    xdi16           : in     std_logic;
    xdi17           : in     std_logic;
    xdi18           : in     std_logic;
    xdi19           : in     std_logic;
    xdi2            : in     std_logic;
    xdi20           : in     std_logic;
    xdi21           : in     std_logic;
    xdi22           : in     std_logic;
    xdi23           : in     std_logic;
    xdi24           : in     std_logic;
    xdi25           : in     std_logic;
    xdi26           : in     std_logic;
    xdi27           : in     std_logic;
    xdi28           : in     std_logic;
    xdi29           : in     std_logic;
    xdi3            : in     std_logic;
    xdi30           : in     std_logic;
    xdi31           : in     std_logic;
    xdi4            : in     std_logic;
    xdi5            : in     std_logic;
    xdi6            : in     std_logic;
    xdi7            : in     std_logic;
    xdi8            : in     std_logic;
    xdi9            : in     std_logic
  );
end entity cadr1_xd;
