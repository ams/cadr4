-- The MIT CADR

library ieee;
use ieee.std_logic_1164.all;

entity cadr4 is
end cadr4;

architecture structural of cadr4 is

begin

  --------------------------------------------------------------------------------

  process
  begin
    wait for 0.1 ns;
  end process;

end structural;
