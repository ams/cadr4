library ieee;
use ieee.std_logic_1164.all;

entity cadr_iram22 is
  port (
    pc0k     : out std_logic;
    pc1k     : out std_logic;
    pc2k     : out std_logic;
    pc3k     : out std_logic;
    pc4k     : out std_logic;
    pc5k     : out std_logic;
    i31      : out std_logic;
    \-iwek\  : in  std_logic;
    \-ice2c\ : in  std_logic;
    iwr31    : in  std_logic;
    pc11k    : out std_logic;
    pc10k    : out std_logic;
    pc9k     : out std_logic;
    pc8k     : out std_logic;
    pc7k     : out std_logic;
    pc6k     : out std_logic;
    i32      : out std_logic;
    iwr32    : in  std_logic;
    i33      : out std_logic;
    iwr33    : in  std_logic;
    i34      : out std_logic;
    iwr34    : in  std_logic;
    i35      : out std_logic;
    iwr35    : in  std_logic;
    i26      : out std_logic;
    iwr26    : in  std_logic;
    i27      : out std_logic;
    iwr27    : in  std_logic;
    i28      : out std_logic;
    iwr28    : in  std_logic;
    i29      : out std_logic;
    iwr29    : in  std_logic;
    i30      : out std_logic;
    iwr30    : in  std_logic;
    \-pcc6\  : in  std_logic;
    \-pcc7\  : in  std_logic;
    \-pcc8\  : in  std_logic;
    \-pcc9\  : in  std_logic;
    \-pcc10\ : in  std_logic;
    \-pcc11\ : in  std_logic;
    \-pcc0\  : in  std_logic;
    \-pcc1\  : in  std_logic;
    \-pcc2\  : in  std_logic;
    \-pcc3\  : in  std_logic;
    \-pcc4\  : in  std_logic;
    \-pcc5\  : in  std_logic;
    i24      : out std_logic;
    iwr24    : in  std_logic;
    i25      : out std_logic;
    iwr25    : in  std_logic
    );
end;
