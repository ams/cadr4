library ieee;
use ieee.std_logic_1164.all;

entity cadr_debug is
  port (
    \-idebug\  : in  std_logic;
    i39        : out std_logic;
    spy7       : in  std_logic;
    spy6       : in  std_logic;
    i38        : out std_logic;
    i37        : out std_logic;
    spy5       : in  std_logic;
    spy4       : in  std_logic;
    i36        : out std_logic;
    \-lddbirh\ : in  std_logic;
    i35        : out std_logic;
    spy3       : in  std_logic;
    spy2       : in  std_logic;
    i34        : out std_logic;
    i33        : out std_logic;
    spy1       : in  std_logic;
    spy0       : in  std_logic;
    i32        : out std_logic;
    i31        : out std_logic;
    spy15      : in  std_logic;
    spy14      : in  std_logic;
    i30        : out std_logic;
    i29        : out std_logic;
    spy13      : in  std_logic;
    spy12      : in  std_logic;
    i28        : out std_logic;
    \-lddbirm\ : in  std_logic;
    i27        : out std_logic;
    spy11      : in  std_logic;
    spy10      : in  std_logic;
    i26        : out std_logic;
    i25        : out std_logic;
    spy9       : in  std_logic;
    spy8       : in  std_logic;
    i24        : out std_logic;
    i23        : out std_logic;
    i22        : out std_logic;
    i21        : out std_logic;
    i20        : out std_logic;
    i19        : out std_logic;
    i18        : out std_logic;
    i17        : out std_logic;
    i16        : out std_logic;
    i15        : out std_logic;
    i14        : out std_logic;
    i13        : out std_logic;
    i12        : out std_logic;
    \-lddbirl\ : in  std_logic;
    i11        : out std_logic;
    i10        : out std_logic;
    i9         : out std_logic;
    i8         : out std_logic;
    i7         : out std_logic;
    i6         : out std_logic;
    i5         : out std_logic;
    i4         : out std_logic;
    i3         : out std_logic;
    i2         : out std_logic;
    i1         : out std_logic;
    i0         : out std_logic;
    i47        : out std_logic;
    i46        : out std_logic;
    i45        : out std_logic;
    i44        : out std_logic;
    i43        : out std_logic;
    i42        : out std_logic;
    i41        : out std_logic;
    i40        : out std_logic);
end;
