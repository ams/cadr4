library ieee;
use ieee.std_logic_1164.all;

entity cadr_bcterm is
  port (
    mem0        : inout std_logic;
    mem1        : inout std_logic;
    mem2        : inout std_logic;
    mem3        : inout std_logic;
    mem4        : inout std_logic;
    mem5        : inout std_logic;
    mem6        : inout std_logic;
    mem7        : inout std_logic;
    mem8        : inout std_logic;
    mem9        : inout std_logic;
    mem10       : inout std_logic;
    mem11       : inout std_logic;
    mem12       : inout std_logic;
    mem13       : inout std_logic;
    mem14       : inout std_logic;
    mem15       : inout std_logic;
    mem16       : inout std_logic;
    mem17       : inout std_logic;
    mem18       : inout std_logic;
    mem19       : inout std_logic;
    mem20       : inout std_logic;
    mem21       : inout std_logic;
    mem22       : inout std_logic;
    mem23       : inout std_logic;
    mem24       : inout std_logic;
    mem25       : inout std_logic;
    mem26       : inout std_logic;
    mem27       : inout std_logic;
    mem28       : inout std_logic;
    mem29       : inout std_logic;
    mem30       : inout std_logic;
    mem31       : inout std_logic;
    \mempar in\ : inout std_logic;
    \-memgrant\ : inout std_logic;
    int         : inout std_logic;
    \-loadmd\   : inout std_logic;
    \-ignpar\   : inout std_logic;
    \-memack\   : inout std_logic);
end;
