library ieee;
use ieee.std_logic_1164.all;

entity cadr_qctl is
  port (
    \-ir0\          : in     std_logic;
    \-ir1\          : in     std_logic;
    \-iralu\        : in     std_logic;
    \-srcq\         : in     std_logic;
    alu31           : in     std_logic;
    q0              : in     std_logic;
    q1              : in     std_logic;
    q10             : in     std_logic;
    q11             : in     std_logic;
    q12             : in     std_logic;
    q13             : in     std_logic;
    q14             : in     std_logic;
    q15             : in     std_logic;
    q16             : in     std_logic;
    q17             : in     std_logic;
    q18             : in     std_logic;
    q19             : in     std_logic;
    q2              : in     std_logic;
    q20             : in     std_logic;
    q21             : in     std_logic;
    q22             : in     std_logic;
    q23             : in     std_logic;
    q24             : in     std_logic;
    q25             : in     std_logic;
    q26             : in     std_logic;
    q27             : in     std_logic;
    q28             : in     std_logic;
    q29             : in     std_logic;
    q3              : in     std_logic;
    q30             : in     std_logic;
    q31             : in     std_logic;
    q4              : in     std_logic;
    q5              : in     std_logic;
    q6              : in     std_logic;
    q7              : in     std_logic;
    q8              : in     std_logic;
    q9              : in     std_logic;
    tse2            : in     std_logic;
    \-alu31\        : out    std_logic;
    \-qdrive\       : out    std_logic;
    mf0             : out    std_logic;
    mf1             : out    std_logic;
    mf10            : out    std_logic;
    mf11            : out    std_logic;
    mf12            : out    std_logic;
    mf13            : out    std_logic;
    mf14            : out    std_logic;
    mf15            : out    std_logic;
    mf16            : out    std_logic;
    mf17            : out    std_logic;
    mf18            : out    std_logic;
    mf19            : out    std_logic;
    mf2             : out    std_logic;
    mf20            : out    std_logic;
    mf21            : out    std_logic;
    mf22            : out    std_logic;
    mf23            : out    std_logic;
    mf24            : out    std_logic;
    mf25            : out    std_logic;
    mf26            : out    std_logic;
    mf27            : out    std_logic;
    mf28            : out    std_logic;
    mf29            : out    std_logic;
    mf3             : out    std_logic;
    mf30            : out    std_logic;
    mf31            : out    std_logic;
    mf4             : out    std_logic;
    mf5             : out    std_logic;
    mf6             : out    std_logic;
    mf7             : out    std_logic;
    mf8             : out    std_logic;
    mf9             : out    std_logic;
    qdrive          : out    std_logic;
    qs0             : out    std_logic;
    qs1             : out    std_logic;
    srcq            : out    std_logic
  );
end entity cadr_qctl;
