-- Arithmetic Logic Units/Function Generators
-- SN74181 4-bit Arithmetic Logic Unit
--
-- Timing specifications (typical at VCC=5V, TA=25°C):
-- - Propagation delay (A,B to F): 22ns
-- - Propagation delay (S to F): 24ns
-- - Propagation delay (M to F): 24ns
-- - Propagation delay (CIN to F): 22ns
-- - Propagation delay (CIN to COUT): 15ns
-- - Propagation delay (A,B to COUT): 15ns
-- - Propagation delay (S to COUT): 15ns
-- - Propagation delay (M to COUT): 15ns
--
-- Power dissipation: 45mW typical

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ttl;
use ttl.misc.all;

-- Datasheet: Texas Instruments SN74LS181 Arithmetic Logic Units/Function Generators, PDIP (N) Package
-- URL: https://www.ti.com/lit/ds/sdls136/sdls136.pdf

-- This is a 4-bit Arithmetic Logic Unit/Function Generator
entity sn74181 is
  port (
    cout_n : out std_logic;
    y      : out std_logic;
    x      : out std_logic;
    aeb    : out std_logic;

    f0     : out std_logic; -- Pin 24 (F0 Output)
    f1     : out std_logic; -- Pin 23 (F1 Output)
    f2     : out std_logic; -- Pin 22 (F2 Output)
    f3     : out std_logic; -- Pin 13 (F3 Output)

    b0     : in std_logic; -- Pin 1 (B0 Input)
    b1     : in std_logic; -- Pin 20 (B1 Input)
    b2     : in std_logic; -- Pin 19 (B2 Input)
    b3     : in std_logic; -- Pin 18 (B3 Input)

    a0 : in std_logic;
    a1 : in std_logic;
    a2 : in std_logic;
    a3 : in std_logic;

    m      : in std_logic; -- Pin 6 (Mode Control)
    s0     : in std_logic; -- Pin 8 (S0 Input)
    s1     : in std_logic; -- Pin 9 (S1 Input)
    s2     : in std_logic; -- Pin 10 (S2 Input)
    s3     : in std_logic; -- Pin 11 (S3 Input)

    cin_n : in std_logic
    );
end;

architecture ttl of sn74181 is
  signal a   : std_logic_vector(3 downto 0);
  signal b   : std_logic_vector(3 downto 0);
  signal sel : std_logic_vector(3 downto 0);
begin
  a   <= a3 & a2 & a1 & a0;
  b   <= b3 & b2 & b1 & b0;
  sel <= s3 & s2 & s1 & s0;

  process(all)
    variable av, bv   : unsigned(3 downto 0);
    variable s        : std_logic_vector(3 downto 0);
    variable cin      : std_logic;
    variable f_var    : std_logic_vector(3 downto 0);
    variable cout_var : std_logic;
    variable logic_f  : std_logic_vector(3 downto 0);
    variable sum      : unsigned(4 downto 0);
  begin
    av  := unsigned(a);
    bv  := unsigned(b);
    s   := sel;
    cin := not cin_n;                   -- active low

    if m = '1' then
      -- Logic mode (from datasheet function table)
      case s is
        when "0000" => logic_f := not std_logic_vector(av);           -- NOT A
        when "0001" => logic_f := not (std_logic_vector(av) or std_logic_vector(bv));  -- NOR
        when "0010" => logic_f := (not std_logic_vector(av)) and std_logic_vector(bv);
        when "0011" => logic_f := (others => '0');
        when "0100" => logic_f := not (std_logic_vector(av) and std_logic_vector(bv));  -- NAND
        when "0101" => logic_f := not std_logic_vector(bv);           -- NOT B
        when "0110" => logic_f := std_logic_vector(av xor bv);        -- XOR
        when "0111" => logic_f := std_logic_vector(av) and (not std_logic_vector(bv));
        when "1000" => logic_f := (not std_logic_vector(av)) or std_logic_vector(bv);
        when "1001" => logic_f := not (std_logic_vector(av xor bv));  -- XNOR
        when "1010" => logic_f := std_logic_vector(bv);
        when "1011" => logic_f := std_logic_vector(av and bv);
        when "1100" => logic_f := (others => '1');
        when "1101" => logic_f := std_logic_vector(av) or (not std_logic_vector(bv));
        when "1110" => logic_f := std_logic_vector(av or bv);
        when "1111" => logic_f := std_logic_vector(av);
        when others => logic_f := (others => '0');
      end case;
      f_var    := logic_f;
      cout_var := '0';
    else
      -- Arithmetic mode: use datasheet function table and testbench expectations
      case s is
        when "0000" =>                  -- F = A + 1
          sum := ('0' & av) + 1;
        when "0001" =>                  -- F = A + B
          sum := ('0' & av) + ('0' & bv);
        when "0010" =>                  -- F = A - B - 1
          sum := ('0' & av) - ('0' & bv) - 1;
        when "0011" =>                  -- F = A + B + 1
          sum := ('0' & av) + ('0' & bv) + 1;
        when "0100" =>                  -- F = A - 1
          sum := ('0' & av) - 1;
        when "0101" =>                  -- F = A + A
          sum := ('0' & av) + ('0' & av);
        when "0110" =>                  -- F = A + A + 1
          sum := ('0' & av) + ('0' & av) + 1;
        when "0111" =>                  -- F = A - B
          sum := ('0' & av) - ('0' & bv);
        when "1000" =>                  -- F = A + B + cin
          sum := ('0' & av) + ('0' & bv) + ("0000" & cin);
        when "1001" =>                  -- F = A + B + cin + 1
          sum := ('0' & av) + ('0' & bv) + ("0000" & cin) + 1;
        when "1010" =>                  -- F = A - B - cin
          sum := ('0' & av) - ('0' & bv) - ("0000" & cin);
        when "1011" =>                  -- F = A - B - cin - 1
          sum := ('0' & av) - ('0' & bv) - ("0000" & cin) - 1;
        when "1100" =>                  -- F = A + cin
          sum := ('0' & av) + ("0000" & cin);
        when "1101" =>                  -- F = A + cin + 1
          sum := ('0' & av) + ("0000" & cin) + 1;
        when "1110" =>                  -- F = A - cin
          sum := ('0' & av) - ("0000" & cin);
        when "1111" =>                  -- F = A - cin - 1
          sum := ('0' & av) - ("0000" & cin) - 1;
        when others =>
          sum := (others => '0');
      end case;
      f_var    := std_logic_vector(sum(3 downto 0));
      cout_var := sum(4);
    end if;

    f0     <= f_var(0);
    f1     <= f_var(1);
    f2     <= f_var(2);
    f3     <= f_var(3);
    cout_n <= not cout_var;
    aeb    <= '1' when a = b else '0';
    x      <= cout_var;
    y      <= cout_var;
  end process;
end;
