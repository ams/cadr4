library ieee;
use ieee.std_logic_1164.all;

-- Dec 14 18:19:44 1980

package cadr_book is

  component cadr_actl is
    port (
      clk3e       : in  std_logic;
      wadr0       : out std_logic;
      ir32        : in  std_logic;
      \-aadr0b\   : out std_logic;
      wadr1       : out std_logic;
      ir33        : in  std_logic;
      \-aadr1b\   : out std_logic;
      \-aadr2b\   : out std_logic;
      ir34        : in  std_logic;
      wadr2       : out std_logic;
      \-aadr3b\   : out std_logic;
      ir35        : in  std_logic;
      wadr3       : out std_logic;
      clk3d       : in  std_logic;
      wadr4       : out std_logic;
      ir36        : in  std_logic;
      \-aadr4b\   : out std_logic;
      wadr5       : out std_logic;
      ir37        : in  std_logic;
      \-aadr5b\   : out std_logic;
      \-aadr6b\   : out std_logic;
      ir38        : in  std_logic;
      wadr6       : out std_logic;
      \-aadr7b\   : out std_logic;
      ir39        : in  std_logic;
      wadr7       : out std_logic;
      \-aadr0a\   : out std_logic;
      \-aadr1a\   : out std_logic;
      \-aadr2a\   : out std_logic;
      \-aadr3a\   : out std_logic;
      \-aadr4a\   : out std_logic;
      \-aadr5a\   : out std_logic;
      \-aadr6a\   : out std_logic;
      \-aadr7a\   : out std_logic;
      wadr8       : out std_logic;
      ir40        : in  std_logic;
      \-aadr8a\   : out std_logic;
      wadr9       : out std_logic;
      ir41        : in  std_logic;
      \-aadr9a\   : out std_logic;
      \-aadr8b\   : out std_logic;
      \-aadr9b\   : out std_logic;
      apass2      : out std_logic;
      \-apass\    : out std_logic;
      tse3a       : in  std_logic;
      \-amemenb\  : out std_logic;
      \-reset\    : in  std_logic;
      ir14        : in  std_logic;
      ir15        : in  std_logic;
      ir16        : in  std_logic;
      ir17        : in  std_logic;
      destmd      : out std_logic;
      destm       : in  std_logic;
      dest        : in  std_logic;
      destd       : out std_logic;
      ir21        : in  std_logic;
      ir20        : in  std_logic;
      ir19        : in  std_logic;
      ir18        : in  std_logic;
      ir23        : in  std_logic;
      ir22        : in  std_logic;
      wp3a        : in  std_logic;
      \-awpa\     : out std_logic;
      \-awpb\     : out std_logic;
      \-awpc\     : out std_logic;
      tse4a       : in  std_logic;
      apassenb    : out std_logic;
      \-apassenb\ : out std_logic;
      apass1      : out std_logic
      );
  end component;

  component cadr_alatch is
    port (
      \-amemenb\  : in  std_logic;
      amem23      : in  std_logic;
      amem22      : in  std_logic;
      a22         : out std_logic;
      a21         : out std_logic;
      amem21      : in  std_logic;
      amem20      : in  std_logic;
      a20         : out std_logic;
      clk3e       : in  std_logic;
      a19         : out std_logic;
      amem19      : in  std_logic;
      amem18      : in  std_logic;
      a18         : out std_logic;
      a17         : out std_logic;
      amem17      : in  std_logic;
      amem16      : in  std_logic;
      a16         : out std_logic;
      \-apassenb\ : in  std_logic;
      l15         : in  std_logic;
      a8          : out std_logic;
      l14         : in  std_logic;
      a9          : out std_logic;
      l13         : in  std_logic;
      a10         : out std_logic;
      l12         : in  std_logic;
      a11         : out std_logic;
      l11         : in  std_logic;
      a12         : out std_logic;
      l10         : in  std_logic;
      a13         : out std_logic;
      l9          : in  std_logic;
      a14         : out std_logic;
      l8          : in  std_logic;
      a15         : out std_logic;
      apassenb    : in  std_logic;
      amem15      : in  std_logic;
      amem14      : in  std_logic;
      amem13      : in  std_logic;
      amem12      : in  std_logic;
      amem11      : in  std_logic;
      amem10      : in  std_logic;
      amem9       : in  std_logic;
      amem8       : in  std_logic;
      l7          : in  std_logic;
      a0          : out std_logic;
      l6          : in  std_logic;
      a1          : out std_logic;
      l5          : in  std_logic;
      a2          : out std_logic;
      l4          : in  std_logic;
      a3          : out std_logic;
      l3          : in  std_logic;
      a4          : out std_logic;
      l2          : in  std_logic;
      a5          : out std_logic;
      l1          : in  std_logic;
      a6          : out std_logic;
      l0          : in  std_logic;
      a7          : out std_logic;
      amem7       : in  std_logic;
      amem6       : in  std_logic;
      amem5       : in  std_logic;
      amem4       : in  std_logic;
      amem3       : in  std_logic;
      amem2       : in  std_logic;
      amem1       : in  std_logic;
      amem0       : in  std_logic;
      a31b        : out std_logic;
      aparity     : out std_logic;
      lparity     : in  std_logic;
      l31         : in  std_logic;
      amemparity  : in  std_logic;
      amem31      : in  std_logic;
      a24         : out std_logic;
      l30         : in  std_logic;
      a25         : out std_logic;
      l29         : in  std_logic;
      a26         : out std_logic;
      l28         : in  std_logic;
      a27         : out std_logic;
      l27         : in  std_logic;
      a28         : out std_logic;
      l26         : in  std_logic;
      a29         : out std_logic;
      l25         : in  std_logic;
      a30         : out std_logic;
      l24         : in  std_logic;
      a31a        : out std_logic;
      amem30      : in  std_logic;
      amem29      : in  std_logic;
      amem28      : in  std_logic;
      amem27      : in  std_logic;
      amem26      : in  std_logic;
      amem25      : in  std_logic;
      amem24      : in  std_logic;
      l23         : in  std_logic;
      l22         : in  std_logic;
      l21         : in  std_logic;
      l20         : in  std_logic;
      l19         : in  std_logic;
      l18         : in  std_logic;
      l17         : in  std_logic;
      l16         : in  std_logic;
      a23         : out std_logic
      );
  end component;

  component cadr_alu0 is
    port (
      a12      : out std_logic;
      m12      : in  std_logic;
      aluf3b   : in  std_logic;
      aluf2b   : in  std_logic;
      aluf1b   : in  std_logic;
      aluf0b   : in  std_logic;
      \-cin12\ : in  std_logic;
      alumode  : in  std_logic;
      alu12    : out std_logic;
      alu13    : out std_logic;
      alu14    : out std_logic;
      alu15    : out std_logic;
      \a=m\    : out std_logic;
      xout15   : out std_logic;
      yout15   : out std_logic;
      a15      : in  std_logic;
      m15      : in  std_logic;
      a14      : in  std_logic;
      m14      : in  std_logic;
      a13      : in  std_logic;
      m13      : in  std_logic;
      a4       : in  std_logic;
      m4       : in  std_logic;
      \-cin4\  : in  std_logic;
      alu4     : out std_logic;
      alu5     : out std_logic;
      alu6     : out std_logic;
      alu7     : out std_logic;
      xout7    : out std_logic;
      yout7    : out std_logic;
      a7       : in  std_logic;
      m7       : in  std_logic;
      a6       : in  std_logic;
      m6       : in  std_logic;
      a5       : in  std_logic;
      m5       : in  std_logic;
      a8       : in  std_logic;
      m8       : in  std_logic;
      \-cin8\  : in  std_logic;
      alu8     : out std_logic;
      alu9     : out std_logic;
      alu10    : out std_logic;
      alu11    : out std_logic;
      xout11   : out std_logic;
      yout11   : out std_logic;
      a11      : in  std_logic;
      m11      : in  std_logic;
      a10      : in  std_logic;
      m10      : in  std_logic;
      a9       : in  std_logic;
      m9       : in  std_logic;
      a0       : in  std_logic;
      m0       : in  std_logic;
      \-cin0\  : in  std_logic;
      alu0     : out std_logic;
      alu1     : out std_logic;
      alu2     : out std_logic;
      alu3     : out std_logic;
      xout3    : out std_logic;
      yout3    : out std_logic;
      a3       : in  std_logic;
      m3       : in  std_logic;
      a2       : in  std_logic;
      m2       : in  std_logic;
      a1       : in  std_logic;
      m1       : in  std_logic
      );
  end component;

  component cadr_alu1 is
    port (
      a31a     : in  std_logic;
      m31b     : out std_logic;
      aluf3a   : in  std_logic;
      aluf2a   : in  std_logic;
      aluf1a   : in  std_logic;
      aluf0a   : in  std_logic;
      \-cin32\ : in  std_logic;
      alumode  : in  std_logic;
      alu32    : out std_logic;
      m31      : in  std_logic;
      a28      : in  std_logic;
      m28      : in  std_logic;
      \-cin28\ : in  std_logic;
      alu28    : out std_logic;
      alu29    : out std_logic;
      alu30    : out std_logic;
      alu31    : out std_logic;
      \a=m\    : out std_logic;
      xout31   : out std_logic;
      yout31   : out std_logic;
      a31b     : in  std_logic;
      a30      : in  std_logic;
      m30      : in  std_logic;
      a29      : in  std_logic;
      m29      : in  std_logic;
      a20      : in  std_logic;
      m20      : in  std_logic;
      \-cin20\ : in  std_logic;
      alu20    : out std_logic;
      alu21    : out std_logic;
      alu22    : out std_logic;
      alu23    : out std_logic;
      xout23   : out std_logic;
      yout23   : out std_logic;
      a23      : in  std_logic;
      m23      : in  std_logic;
      a22      : in  std_logic;
      m22      : in  std_logic;
      a21      : in  std_logic;
      m21      : in  std_logic;
      a24      : in  std_logic;
      m24      : in  std_logic;
      \-cin24\ : in  std_logic;
      alu24    : out std_logic;
      alu25    : out std_logic;
      alu26    : out std_logic;
      alu27    : out std_logic;
      xout27   : out std_logic;
      yout27   : out std_logic;
      a27      : in  std_logic;
      m27      : in  std_logic;
      a26      : in  std_logic;
      m26      : in  std_logic;
      a25      : in  std_logic;
      m25      : in  std_logic;
      a16      : in  std_logic;
      m16      : in  std_logic;
      \-cin16\ : in  std_logic;
      alu16    : out std_logic;
      alu17    : out std_logic;
      alu18    : out std_logic;
      alu19    : out std_logic;
      xout19   : out std_logic;
      yout19   : out std_logic;
      a19      : in  std_logic;
      m19      : in  std_logic;
      a18      : in  std_logic;
      m18      : in  std_logic;
      a17      : in  std_logic;
      m17      : in  std_logic
      );
  end component;

  component cadr_aluc4 is
    port (
      \-aluf0\          : out std_logic;
      aluf0b            : out std_logic;
      \-aluf1\          : out std_logic;
      aluf1b            : out std_logic;
      aluf2b            : out std_logic;
      \-aluf2\          : out std_logic;
      aluf3b            : out std_logic;
      \-aluf3\          : out std_logic;
      aluf0a            : out std_logic;
      aluf1a            : out std_logic;
      aluf2a            : out std_logic;
      aluf3a            : out std_logic;
      yy1               : out std_logic;
      xx1               : out std_logic;
      yy0               : out std_logic;
      xx0               : out std_logic;
      \-cin32\          : out std_logic;
      \-cin16\          : out std_logic;
      \-cin0\           : out std_logic;
      yout23            : in  std_logic;
      xout23            : in  std_logic;
      yout19            : in  std_logic;
      xout19            : in  std_logic;
      yout31            : out std_logic;
      xout31            : out std_logic;
      \-cin28\          : out std_logic;
      \-cin24\          : out std_logic;
      \-cin20\          : out std_logic;
      yout27            : in  std_logic;
      xout27            : in  std_logic;
      yout7             : in  std_logic;
      xout7             : in  std_logic;
      yout3             : in  std_logic;
      xout3             : in  std_logic;
      yout15            : out std_logic;
      xout15            : out std_logic;
      \-cin12\          : out std_logic;
      \-cin8\           : out std_logic;
      \-cin4\           : out std_logic;
      yout11            : in  std_logic;
      xout11            : in  std_logic;
      alusub            : out std_logic;
      \-ir3\            : out std_logic;
      \-ir4\            : out std_logic;
      aluadd            : out std_logic;
      ir6               : in  std_logic;
      ir5               : in  std_logic;
      ir7               : in  std_logic;
      \-alumode\        : out std_logic;
      \-ir2\            : out std_logic;
      irjump            : in  std_logic;
      alumode           : out std_logic;
      \-divposlasttime\ : out std_logic;
      q0                : in  std_logic;
      \-div\            : in  std_logic;
      divsubcond        : out std_logic;
      divaddcond        : out std_logic;
      a31b              : in  std_logic;
      \-a31\            : out std_logic;
      ir4               : in  std_logic;
      ir3               : in  std_logic;
      ir2               : in  std_logic;
      \-ir1\            : out std_logic;
      ir1               : in  std_logic;
      \-ir0\            : out std_logic;
      ir0               : in  std_logic;
      a31a              : in  std_logic;
      \-mulnop\         : out std_logic;
      \-irjump\         : in  std_logic;
      \-mul\            : in  std_logic;
      osel1a            : out std_logic;
      \-ir13\           : in  std_logic;
      \-iralu\          : in  std_logic;
      osel0a            : out std_logic;
      \-ir12\           : in  std_logic;
      osel1b            : out std_logic;
      osel0b            : out std_logic
      );
  end component;

  component cadr_amem0 is
    port (
      \-aadr0b\  : in  std_logic;
      \-aadr1b\  : in  std_logic;
      \-aadr2b\  : in  std_logic;
      \-aadr3b\  : in  std_logic;
      \-aadr4b\  : in  std_logic;
      amem22     : out std_logic;
      \-aadr5b\  : in  std_logic;
      \-aadr6b\  : in  std_logic;
      \-aadr7b\  : in  std_logic;
      \-aadr8b\  : in  std_logic;
      \-aadr9b\  : in  std_logic;
      \-awpa\    : in  std_logic;
      l22        : in  std_logic;
      amem20     : out std_logic;
      \-awpb\    : in  std_logic;
      l20        : in  std_logic;
      amem18     : out std_logic;
      l18        : in  std_logic;
      amem16     : out std_logic;
      l16        : in  std_logic;
      amem23     : out std_logic;
      l23        : in  std_logic;
      amem21     : out std_logic;
      l21        : in  std_logic;
      amem19     : out std_logic;
      l19        : in  std_logic;
      amem17     : out std_logic;
      l17        : in  std_logic;
      amemparity : out std_logic;
      lparity    : in  std_logic;
      amem30     : out std_logic;
      l30        : in  std_logic;
      amem28     : out std_logic;
      l28        : in  std_logic;
      amem26     : out std_logic;
      l26        : in  std_logic;
      amem24     : out std_logic;
      l24        : in  std_logic;
      amem31     : out std_logic;
      l31        : in  std_logic;
      amem29     : out std_logic;
      l29        : in  std_logic;
      amem27     : out std_logic;
      l27        : in  std_logic;
      amem25     : out std_logic;
      l25        : in  std_logic
      );
  end component;

  component cadr_amem1 is
    port (
      \-aadr0a\ : in  std_logic;
      \-aadr1a\ : in  std_logic;
      \-aadr2a\ : in  std_logic;
      \-aadr3a\ : in  std_logic;
      \-aadr4a\ : in  std_logic;
      amem6     : out std_logic;
      \-aadr5a\ : in  std_logic;
      \-aadr6a\ : in  std_logic;
      \-aadr7a\ : in  std_logic;
      \-aadr8a\ : in  std_logic;
      \-aadr9a\ : in  std_logic;
      \-awpc\   : in  std_logic;
      l6        : in  std_logic;
      amem4     : out std_logic;
      l4        : in  std_logic;
      amem2     : out std_logic;
      l2        : in  std_logic;
      amem0     : out std_logic;
      l0        : in  std_logic;
      amem7     : out std_logic;
      l7        : in  std_logic;
      amem5     : out std_logic;
      l5        : in  std_logic;
      amem3     : out std_logic;
      l3        : in  std_logic;
      amem1     : out std_logic;
      l1        : in  std_logic;
      amem14    : out std_logic;
      \-awpb\   : in  std_logic;
      l14       : in  std_logic;
      amem12    : out std_logic;
      l12       : in  std_logic;
      amem10    : out std_logic;
      l10       : in  std_logic;
      amem8     : out std_logic;
      l8        : in  std_logic;
      amem15    : out std_logic;
      l15       : in  std_logic;
      amem13    : out std_logic;
      l13       : in  std_logic;
      amem11    : out std_logic;
      l11       : in  std_logic;
      amem9     : out std_logic;
      l9        : in  std_logic
      );
  end component;

  component cadr_apar is
    port (
      a26       : in  std_logic;
      a27       : in  std_logic;
      a28       : in  std_logic;
      a29       : in  std_logic;
      a30       : in  std_logic;
      a31b      : in  std_logic;
      aparity   : in  std_logic;
      aparok    : out std_logic;
      aparl     : out std_logic;
      aparm     : out std_logic;
      a24       : in  std_logic;
      a25       : in  std_logic;
      a17       : in  std_logic;
      a18       : in  std_logic;
      a19       : in  std_logic;
      a20       : in  std_logic;
      a21       : in  std_logic;
      a22       : in  std_logic;
      a23       : in  std_logic;
      a12       : in  std_logic;
      a13       : in  std_logic;
      a14       : in  std_logic;
      a15       : in  std_logic;
      a16       : in  std_logic;
      a5        : in  std_logic;
      a6        : in  std_logic;
      a7        : in  std_logic;
      a8        : in  std_logic;
      a9        : in  std_logic;
      a10       : in  std_logic;
      a11       : in  std_logic;
      a0        : in  std_logic;
      a1        : in  std_logic;
      a2        : in  std_logic;
      a3        : in  std_logic;
      a4        : in  std_logic;
      m17       : in  std_logic;
      m18       : in  std_logic;
      m19       : in  std_logic;
      m20       : in  std_logic;
      m21       : in  std_logic;
      m22       : in  std_logic;
      m23       : in  std_logic;
      mparm     : out std_logic;
      m12       : in  std_logic;
      m13       : in  std_logic;
      m14       : in  std_logic;
      m15       : in  std_logic;
      m16       : in  std_logic;
      m5        : in  std_logic;
      m6        : in  std_logic;
      m7        : in  std_logic;
      m8        : in  std_logic;
      m9        : in  std_logic;
      m10       : in  std_logic;
      m11       : in  std_logic;
      mparl     : out std_logic;
      m0        : in  std_logic;
      m1        : in  std_logic;
      m2        : in  std_logic;
      m3        : in  std_logic;
      m4        : in  std_logic;
      mpareven  : out std_logic;
      srcm      : in  std_logic;
      mmemparok : out std_logic;
      pdlenb    : in  std_logic;
      pdlparok  : out std_logic;
      m26       : in  std_logic;
      m27       : in  std_logic;
      m28       : in  std_logic;
      m29       : in  std_logic;
      m30       : in  std_logic;
      m31       : in  std_logic;
      mparity   : in  std_logic;
      mparodd   : out std_logic;
      m24       : in  std_logic;
      m25       : in  std_logic
      );
  end component;

-- component cadr_bcpins is
-- end component;

  component cadr_bcterm is
    port (
      mem0        : out std_logic;
      mem1        : out std_logic;
      mem2        : out std_logic;
      mem3        : out std_logic;
      mem4        : out std_logic;
      mem5        : out std_logic;
      mem6        : out std_logic;
      mem7        : out std_logic;
      mem8        : out std_logic;
      mem9        : out std_logic;
      mem10       : out std_logic;
      mem11       : out std_logic;
      mem12       : out std_logic;
      mem13       : out std_logic;
      mem14       : out std_logic;
      mem15       : out std_logic;
      mem16       : out std_logic;
      mem17       : out std_logic;
      mem18       : out std_logic;
      mem19       : out std_logic;
      mem20       : out std_logic;
      mem21       : out std_logic;
      mem22       : out std_logic;
      mem23       : out std_logic;
      mem24       : out std_logic;
      mem25       : out std_logic;
      mem26       : out std_logic;
      mem27       : out std_logic;
      mem28       : out std_logic;
      mem29       : out std_logic;
      mem30       : out std_logic;
      mem31       : out std_logic;
      \mempar in\ : out std_logic;
      \-memgrant\ : out std_logic;
      int         : out std_logic;
      \-loadmd\   : out std_logic;
      \-ignpar\   : out std_logic;
      \-memack\   : out std_logic
      );
  end component;

-- component cadr_caps is
-- end component;

  component cadr_clockd is
    port (
      \-clk1\        : out std_logic;
      clk1a          : out std_logic;
      reset          : in  std_logic;
      \-reset\       : out std_logic;
      mclk1a         : out std_logic;
      \-mclk1\       : out std_logic;
      mclk1          : in  std_logic;
      clk1           : in  std_logic;
      \-wp1\         : in  std_logic;
      wp1b           : out std_logic;
      wp1a           : out std_logic;
      tse1b          : out std_logic;
      \-tse1\        : in  std_logic;
      tse1a          : out std_logic;
      \-upperhighok\ : out std_logic;
      lcry3          : in  std_logic;
      \-lcry3\       : out std_logic;
      clk2           : in  std_logic;
      \-clk2c\       : out std_logic;
      \-clk2a\       : out std_logic;
      wp2            : out std_logic;
      \-wp2\         : in  std_logic;
      tse2           : out std_logic;
      \-tse2\        : in  std_logic;
      clk2a          : out std_logic;
      clk2b          : out std_logic;
      clk2c          : out std_logic;
      \-clk3a\       : out std_logic;
      clk3a          : out std_logic;
      clk3b          : out std_logic;
      clk3c          : out std_logic;
      clk3           : in  std_logic;
      \-clk3g\       : out std_logic;
      \-clk3d\       : out std_logic;
      wp3a           : out std_logic;
      \-wp3\         : in  std_logic;
      tse3a          : out std_logic;
      \-tse3\        : in  std_logic;
      clk3d          : out std_logic;
      clk3e          : out std_logic;
      clk3f          : out std_logic;
      \-clk4a\       : out std_logic;
      clk4a          : out std_logic;
      clk4b          : out std_logic;
      clk4c          : out std_logic;
      clk4           : in  std_logic;
      \-clk4e\       : out std_logic;
      \-clk4d\       : out std_logic;
      wp4c           : out std_logic;
      \-wp4\         : in  std_logic;
      wp4b           : out std_logic;
      wp4a           : out std_logic;
      clk4d          : out std_logic;
      clk4e          : out std_logic;
      clk4f          : out std_logic;
      \-tse4\        : in  std_logic;
      tse4b          : out std_logic;
      tse4a          : out std_logic;
      srcpdlptr      : out std_logic;
      \-srcpdlptr\   : in  std_logic;
      srcpdlidx      : out std_logic;
      \-srcpdlidx\   : in  std_logic
      );
  end component;

  component cadr_contrl is
    port (
      spushd           : out std_logic;
      tse3a            : in  std_logic;
      spcwpass         : out std_logic;
      \-ipopj\         : out std_logic;
      \-iwrited\       : out std_logic;
      \-popj\          : out std_logic;
      spcdrive         : out std_logic;
      spcenb           : out std_logic;
      \-reset\         : in  std_logic;
      inop             : out std_logic;
      \-inop\          : out std_logic;
      n                : out std_logic;
      clk3c            : in  std_logic;
      \-spushd\        : out std_logic;
      spush            : out std_logic;
      iwrite           : out std_logic;
      iwrited          : out std_logic;
      \-srcspc\        : in  std_logic;
      \-srcspcpop\     : in  std_logic;
      \-spcdrive\      : out std_logic;
      \-spcpass\       : out std_logic;
      \-spcwpass\      : out std_logic;
      ir42             : in  std_logic;
      \-nop\           : out std_logic;
      nop              : out std_logic;
      \-srcspcpopreal\ : out std_logic;
      \-nopa\          : out std_logic;
      \-nop11\         : in  std_logic;
      \-irdisp\        : in  std_logic;
      dr               : in  std_logic;
      \-ignpopj\       : out std_logic;
      \-destspc\       : out std_logic;
      destspc          : out std_logic;
      dp               : in  std_logic;
      \-dfall\         : out std_logic;
      \-trap\          : in  std_logic;
      irdisp           : in  std_logic;
      \-funct2\        : in  std_logic;
      dispenb          : out std_logic;
      irjump           : in  std_logic;
      ir6              : in  std_logic;
      jfalse           : out std_logic;
      jcalf            : out std_logic;
      ir8              : in  std_logic;
      jretf            : out std_logic;
      jret             : out std_logic;
      ir7              : in  std_logic;
      dn               : out std_logic;
      \-jcond\         : in  std_logic;
      jcond            : in  std_logic;
      \-ir6\           : out std_logic;
      \-dr\            : out std_logic;
      \-spush\         : out std_logic;
      pcs1             : out std_logic;
      popj             : out std_logic;
      \-dp\            : out std_logic;
      \-spop\          : out std_logic;
      \-ir8\           : out std_logic;
      ir9              : in  std_logic;
      pcs0             : out std_logic;
      \-spcnt\         : out std_logic;
      \-destspcd\      : out std_logic;
      destspcd         : out std_logic;
      \-swpb\          : out std_logic;
      \-swpa\          : out std_logic;
      wp4c             : in  std_logic
      );
  end component;

-- component cadr_cpins is
-- end component;

  component cadr_dram0 is
    port (
      wp2         : in  std_logic;
      dispwr      : in  std_logic;
      \-dwea\     : out std_logic;
      \-dadr10a\  : out std_logic;
      dadr10a     : out std_logic;
      ir22b       : in  std_logic;
      \-dadr9a\   : out std_logic;
      ir21b       : in  std_logic;
      \-dadr8a\   : out std_logic;
      ir20b       : in  std_logic;
      \-dadr7a\   : out std_logic;
      ir19b       : out std_logic;
      ir12b       : out std_logic;
      vmo19       : in  std_logic;
      ir9b        : in  std_logic;
      r0          : in  std_logic;
      dmask0      : in  std_logic;
      \-dmapbenb\ : in  std_logic;
      \-dadr0a\   : out std_logic;
      vmo18       : in  std_logic;
      ir8b        : in  std_logic;
      ir12        : in  std_logic;
      ir13        : in  std_logic;
      ir18b       : out std_logic;
      ir14        : in  std_logic;
      ir17b       : out std_logic;
      ir15        : in  std_logic;
      ir16b       : out std_logic;
      ir16        : in  std_logic;
      ir15b       : out std_logic;
      ir17        : in  std_logic;
      ir14b       : out std_logic;
      ir18        : in  std_logic;
      ir13b       : out std_logic;
      ir19        : in  std_logic;
      \-dadr1a\   : out std_logic;
      \-dadr2a\   : out std_logic;
      \-dadr3a\   : out std_logic;
      \-dadr4a\   : out std_logic;
      dpc5        : out std_logic;
      \-dadr5a\   : out std_logic;
      \-dadr6a\   : out std_logic;
      aa5         : in  std_logic;
      dpc4        : out std_logic;
      aa4         : in  std_logic;
      r3          : in  std_logic;
      dmask6      : in  std_logic;
      r6          : in  std_logic;
      dmask3      : in  std_logic;
      dpc3        : out std_logic;
      aa3         : in  std_logic;
      dpc2        : out std_logic;
      aa2         : in  std_logic;
      r2          : in  std_logic;
      dmask5      : in  std_logic;
      r5          : in  std_logic;
      dmask2      : in  std_logic;
      dpc1        : out std_logic;
      aa1         : in  std_logic;
      dpc0        : out std_logic;
      aa0         : in  std_logic;
      r1          : in  std_logic;
      dmask4      : in  std_logic;
      r4          : in  std_logic;
      dmask1      : in  std_logic
      );
  end component;

  component cadr_dram1 is
    port (
      wp2         : in  std_logic;
      dispwr      : in  std_logic;
      \-dweb\     : out std_logic;
      \-vmo19\    : out std_logic;
      vmo19       : out std_logic;
      \-vmo18\    : out std_logic;
      vmo18       : out std_logic;
      \-dadr9b\   : out std_logic;
      ir21b       : out std_logic;
      \-dadr8b\   : out std_logic;
      ir20b       : out std_logic;
      \-dadr7b\   : out std_logic;
      ir19b       : in  std_logic;
      ir12b       : in  std_logic;
      ir9b        : out std_logic;
      r0          : in  std_logic;
      dmask0      : in  std_logic;
      \-dmapbenb\ : in  std_logic;
      \-dadr0b\   : out std_logic;
      ir8b        : out std_logic;
      dadr10a     : in  std_logic;
      \-dadr1b\   : out std_logic;
      \-dadr2b\   : out std_logic;
      \-dadr3b\   : out std_logic;
      \-dadr4b\   : out std_logic;
      dpc11       : out std_logic;
      \-dadr5b\   : out std_logic;
      \-dadr6b\   : out std_logic;
      aa11        : in  std_logic;
      \-dadr10a\  : in  std_logic;
      dpc10       : out std_logic;
      aa10        : in  std_logic;
      r3          : in  std_logic;
      ir18b       : in  std_logic;
      dmask6      : in  std_logic;
      r6          : in  std_logic;
      ir15b       : in  std_logic;
      dmask3      : in  std_logic;
      dpc9        : out std_logic;
      aa9         : in  std_logic;
      dadr10c     : in  std_logic;
      dpc8        : out std_logic;
      aa8         : in  std_logic;
      \-dadr10c\  : in  std_logic;
      r2          : in  std_logic;
      ir17b       : in  std_logic;
      dmask5      : in  std_logic;
      r5          : in  std_logic;
      ir14b       : in  std_logic;
      dmask2      : in  std_logic;
      dpc7        : out std_logic;
      aa7         : in  std_logic;
      dpc6        : out std_logic;
      aa6         : in  std_logic;
      r1          : in  std_logic;
      ir16b       : in  std_logic;
      dmask4      : in  std_logic;
      r4          : in  std_logic;
      ir13b       : in  std_logic;
      dmask1      : in  std_logic;
      ir20        : in  std_logic;
      ir21        : in  std_logic;
      ir22        : in  std_logic;
      ir8         : in  std_logic;
      ir9         : in  std_logic;
      ir22b       : out std_logic
      );
  end component;

  component cadr_dram2 is
    port (
      dadr10c     : out std_logic;
      \-dadr0c\   : out std_logic;
      \-dadr1c\   : out std_logic;
      \-dadr2c\   : out std_logic;
      \-dadr3c\   : out std_logic;
      \-dadr4c\   : out std_logic;
      dpar        : out std_logic;
      \-dadr5c\   : out std_logic;
      \-dadr6c\   : out std_logic;
      \-dadr7c\   : out std_logic;
      \-dadr8c\   : out std_logic;
      \-dadr9c\   : out std_logic;
      \-dwec\     : out std_logic;
      aa17        : in  std_logic;
      \-dadr10c\  : out std_logic;
      dr          : out std_logic;
      aa16        : in  std_logic;
      r3          : in  std_logic;
      ir18b       : in  std_logic;
      dmask6      : in  std_logic;
      r6          : in  std_logic;
      ir15b       : in  std_logic;
      dmask3      : in  std_logic;
      dp          : out std_logic;
      aa15        : in  std_logic;
      dn          : out std_logic;
      aa14        : in  std_logic;
      r2          : in  std_logic;
      ir17b       : in  std_logic;
      dmask5      : in  std_logic;
      r5          : in  std_logic;
      ir14b       : in  std_logic;
      dmask2      : in  std_logic;
      dpc13       : out std_logic;
      aa13        : in  std_logic;
      dpc12       : out std_logic;
      aa12        : in  std_logic;
      r1          : in  std_logic;
      ir16b       : in  std_logic;
      dmask4      : in  std_logic;
      r4          : in  std_logic;
      ir13b       : in  std_logic;
      dmask1      : in  std_logic;
      ir12b       : in  std_logic;
      vmo19       : in  std_logic;
      ir9b        : in  std_logic;
      r0          : in  std_logic;
      dmask0      : in  std_logic;
      \-dmapbenb\ : in  std_logic;
      vmo18       : in  std_logic;
      ir8b        : in  std_logic;
      ir22b       : in  std_logic;
      ir21b       : in  std_logic;
      ir20b       : in  std_logic;
      ir19b       : in  std_logic;
      dispwr      : in  std_logic;
      wp2         : in  std_logic
      );
  end component;

  component cadr_dspctl is
    port (
      dmask0      : out std_logic;
      dmask1      : out std_logic;
      dmask2      : out std_logic;
      dmask3      : out std_logic;
      dmask4      : out std_logic;
      dmask5      : out std_logic;
      dmask6      : out std_logic;
      ir5         : in  std_logic;
      ir6         : in  std_logic;
      ir7         : in  std_logic;
      \-irdisp\   : in  std_logic;
      dc6         : out std_logic;
      ir38        : in  std_logic;
      ir39        : in  std_logic;
      dc7         : out std_logic;
      ir40        : in  std_logic;
      dc8         : out std_logic;
      clk3e       : in  std_logic;
      dc9         : out std_logic;
      ir41        : in  std_logic;
      dc0         : out std_logic;
      ir32        : in  std_logic;
      ir33        : in  std_logic;
      dc1         : out std_logic;
      ir34        : in  std_logic;
      dc2         : out std_logic;
      dc3         : out std_logic;
      ir35        : in  std_logic;
      dc4         : out std_logic;
      ir36        : in  std_logic;
      ir37        : in  std_logic;
      dc5         : out std_logic;
      dpareven    : out std_logic;
      dispenb     : in  std_logic;
      dparok      : out std_logic;
      \-dparh\    : out std_logic;
      dparl       : out std_logic;
      aa16        : out std_logic;
      aa17        : out std_logic;
      a17         : in  std_logic;
      a16         : in  std_logic;
      a15         : in  std_logic;
      aa8         : out std_logic;
      a14         : in  std_logic;
      aa9         : out std_logic;
      a13         : in  std_logic;
      aa10        : out std_logic;
      a12         : in  std_logic;
      aa11        : out std_logic;
      a11         : in  std_logic;
      aa12        : out std_logic;
      a10         : in  std_logic;
      aa13        : out std_logic;
      a9          : in  std_logic;
      aa14        : out std_logic;
      a8          : in  std_logic;
      aa15        : out std_logic;
      a7          : in  std_logic;
      aa0         : out std_logic;
      a6          : in  std_logic;
      aa1         : out std_logic;
      a5          : in  std_logic;
      aa2         : out std_logic;
      a4          : in  std_logic;
      aa3         : out std_logic;
      a3          : in  std_logic;
      aa4         : out std_logic;
      a2          : in  std_logic;
      aa5         : out std_logic;
      a1          : in  std_logic;
      aa6         : out std_logic;
      a0          : in  std_logic;
      aa7         : out std_logic;
      \-dmapbenb\ : out std_logic;
      ir8         : in  std_logic;
      ir9         : in  std_logic;
      dispwr      : out std_logic;
      \-funct2\   : in  std_logic;
      dpc9        : in  std_logic;
      dpc10       : in  std_logic;
      dpc11       : in  std_logic;
      dpc12       : in  std_logic;
      dpc13       : in  std_logic;
      dn          : in  std_logic;
      dp          : in  std_logic;
      dr          : in  std_logic;
      dpar        : in  std_logic;
      dpc0        : in  std_logic;
      dpc1        : in  std_logic;
      dpc2        : in  std_logic;
      dpc3        : in  std_logic;
      dpc4        : in  std_logic;
      dpc5        : in  std_logic;
      dpc6        : in  std_logic;
      dpc7        : in  std_logic;
      dpc8        : in  std_logic
      );
  end component;

  component cadr_flag is
    port (
      ir45                : in  std_logic;
      \-nopa\             : in  std_logic;
      \-ilong\            : out std_logic;
      ob29                : in  std_logic;
      \lc byte mode\      : out std_logic;
      ob28                : in  std_logic;
      \prog.unibus.reset\ : out std_logic;
      clk3c               : in  std_logic;
      \int.enable\        : out std_logic;
      ob27                : in  std_logic;
      \sequence.break\    : out std_logic;
      ob26                : in  std_logic;
      \-destintctl\       : in  std_logic;
      \-reset\            : in  std_logic;
      \-statbit\          : out std_logic;
      ir46                : in  std_logic;
      \a=m\               : in  std_logic;
      alu32               : in  std_logic;
      aluneg              : out std_logic;
      r0                  : in  std_logic;
      jcond               : out std_logic;
      \-jcond\            : out std_logic;
      conds2              : out std_logic;
      conds1              : out std_logic;
      conds0              : out std_logic;
      \pgf.or.int.or.sb\  : out std_logic;
      \pgf.or.int\        : out std_logic;
      \-vmaok\            : in  std_logic;
      ir2                 : in  std_logic;
      ir5                 : in  std_logic;
      ir1                 : in  std_logic;
      ir0                 : in  std_logic;
      \-alu32\            : out std_logic;
      sint                : out std_logic;
      sintr               : in  std_logic
      );
  end component;

  component cadr_ior is
    port (
      i12   : in  std_logic;
      ob12  : in  std_logic;
      iob12 : out std_logic;
      i13   : in  std_logic;
      ob13  : in  std_logic;
      iob13 : out std_logic;
      iob14 : out std_logic;
      i14   : in  std_logic;
      ob14  : in  std_logic;
      iob15 : out std_logic;
      i15   : in  std_logic;
      ob15  : in  std_logic;
      i8    : in  std_logic;
      ob8   : in  std_logic;
      iob8  : out std_logic;
      i9    : in  std_logic;
      ob9   : in  std_logic;
      iob9  : out std_logic;
      iob10 : out std_logic;
      i10   : in  std_logic;
      ob10  : in  std_logic;
      iob11 : out std_logic;
      i11   : in  std_logic;
      ob11  : in  std_logic;
      i4    : in  std_logic;
      ob4   : in  std_logic;
      iob4  : out std_logic;
      i5    : in  std_logic;
      ob5   : in  std_logic;
      iob5  : out std_logic;
      iob6  : out std_logic;
      i6    : in  std_logic;
      ob6   : in  std_logic;
      iob7  : out std_logic;
      i7    : in  std_logic;
      ob7   : in  std_logic;
      i0    : in  std_logic;
      ob0   : in  std_logic;
      iob0  : out std_logic;
      i1    : in  std_logic;
      iob1  : out std_logic;
      iob2  : out std_logic;
      i2    : in  std_logic;
      ob2   : in  std_logic;
      iob3  : out std_logic;
      i3    : in  std_logic;
      ob3   : in  std_logic;
      i20   : in  std_logic;
      ob20  : in  std_logic;
      iob20 : out std_logic;
      i21   : in  std_logic;
      ob21  : in  std_logic;
      iob21 : out std_logic;
      iob22 : out std_logic;
      i22   : in  std_logic;
      ob22  : in  std_logic;
      iob23 : out std_logic;
      i23   : in  std_logic;
      ob23  : in  std_logic;
      i16   : in  std_logic;
      ob16  : in  std_logic;
      iob16 : out std_logic;
      i17   : in  std_logic;
      ob17  : in  std_logic;
      iob17 : out std_logic;
      iob18 : out std_logic;
      i18   : in  std_logic;
      ob18  : in  std_logic;
      iob19 : out std_logic;
      i19   : in  std_logic;
      ob19  : in  std_logic;
      i44   : in  std_logic;
      iob44 : out std_logic;
      i45   : in  std_logic;
      iob45 : out std_logic;
      iob46 : out std_logic;
      i46   : in  std_logic;
      iob47 : out std_logic;
      i47   : in  std_logic;
      i40   : in  std_logic;
      iob40 : out std_logic;
      i41   : in  std_logic;
      iob41 : out std_logic;
      iob42 : out std_logic;
      i42   : in  std_logic;
      iob43 : out std_logic;
      i43   : in  std_logic;
      i36   : in  std_logic;
      iob36 : out std_logic;
      i37   : in  std_logic;
      iob37 : out std_logic;
      iob38 : out std_logic;
      i38   : in  std_logic;
      iob39 : out std_logic;
      i39   : in  std_logic;
      i32   : in  std_logic;
      iob32 : out std_logic;
      i33   : in  std_logic;
      iob33 : out std_logic;
      iob34 : out std_logic;
      i34   : in  std_logic;
      iob35 : out std_logic;
      i35   : in  std_logic;
      i28   : in  std_logic;
      iob28 : out std_logic;
      i29   : in  std_logic;
      iob29 : out std_logic;
      iob30 : out std_logic;
      i30   : in  std_logic;
      iob31 : out std_logic;
      i31   : in  std_logic;
      i24   : in  std_logic;
      ob24  : in  std_logic;
      iob24 : out std_logic;
      i25   : in  std_logic;
      ob25  : in  std_logic;
      iob25 : out std_logic;
      iob26 : out std_logic;
      i26   : in  std_logic;
      iob27 : out std_logic;
      i27   : in  std_logic;
      ob1   : in  std_logic
      );
  end component;

  component cadr_ipar is
    port (
      ir41    : in  std_logic;
      ir42    : in  std_logic;
      ir43    : in  std_logic;
      ir44    : in  std_logic;
      ir45    : in  std_logic;
      ir46    : in  std_logic;
      ir47    : in  std_logic;
      ipar3   : out std_logic;
      ir36    : in  std_logic;
      ir37    : in  std_logic;
      ir38    : in  std_logic;
      ir39    : in  std_logic;
      ir40    : in  std_logic;
      ir5     : in  std_logic;
      ir6     : in  std_logic;
      ir7     : in  std_logic;
      ir8     : in  std_logic;
      ir9     : in  std_logic;
      ir10    : in  std_logic;
      ir11    : in  std_logic;
      ipar0   : out std_logic;
      ir0     : in  std_logic;
      ir1     : in  std_logic;
      ir2     : in  std_logic;
      ir3     : in  std_logic;
      ir4     : in  std_logic;
      ir29    : in  std_logic;
      ir30    : in  std_logic;
      ir31    : in  std_logic;
      ir32    : in  std_logic;
      ir33    : in  std_logic;
      ir34    : in  std_logic;
      ir35    : in  std_logic;
      ipar2   : out std_logic;
      ir24    : in  std_logic;
      ir25    : in  std_logic;
      ir26    : in  std_logic;
      ir27    : in  std_logic;
      ir28    : in  std_logic;
      iparity : out std_logic;
      ipar1   : out std_logic;
      ir48    : in  std_logic;
      ir17    : in  std_logic;
      ir18    : in  std_logic;
      ir19    : in  std_logic;
      ir20    : in  std_logic;
      ir21    : in  std_logic;
      ir22    : in  std_logic;
      ir23    : in  std_logic;
      ir12    : in  std_logic;
      ir13    : in  std_logic;
      ir14    : in  std_logic;
      ir15    : in  std_logic;
      ir16    : in  std_logic;
      imodd   : in  std_logic;
      iparok  : out std_logic
      );
  end component;

  component cadr_ireg is
    port (
      \-destimod0\ : in  std_logic;
      ir15         : out std_logic;
      iob15        : in  std_logic;
      i15          : in  std_logic;
      i14          : in  std_logic;
      iob14        : in  std_logic;
      ir14         : out std_logic;
      clk3a        : in  std_logic;
      ir13         : out std_logic;
      iob13        : in  std_logic;
      i13          : in  std_logic;
      i12          : in  std_logic;
      iob12        : in  std_logic;
      ir12         : out std_logic;
      ir11         : out std_logic;
      iob11        : in  std_logic;
      i11          : in  std_logic;
      i10          : in  std_logic;
      iob10        : in  std_logic;
      ir10         : out std_logic;
      ir9          : out std_logic;
      iob9         : in  std_logic;
      i9           : in  std_logic;
      i8           : in  std_logic;
      iob8         : in  std_logic;
      ir8          : out std_logic;
      ir7          : out std_logic;
      iob7         : in  std_logic;
      i7           : in  std_logic;
      i6           : in  std_logic;
      iob6         : in  std_logic;
      ir6          : out std_logic;
      ir5          : out std_logic;
      iob5         : in  std_logic;
      i5           : in  std_logic;
      i4           : in  std_logic;
      iob4         : in  std_logic;
      ir4          : out std_logic;
      ir3          : out std_logic;
      iob3         : in  std_logic;
      i3           : in  std_logic;
      i2           : in  std_logic;
      iob2         : in  std_logic;
      ir2          : out std_logic;
      ir1          : out std_logic;
      iob1         : in  std_logic;
      i1           : in  std_logic;
      i0           : in  std_logic;
      iob0         : in  std_logic;
      ir0          : out std_logic;
      ir23         : out std_logic;
      iob23        : in  std_logic;
      i23          : in  std_logic;
      i22          : in  std_logic;
      iob22        : in  std_logic;
      ir22         : out std_logic;
      clk3b        : in  std_logic;
      ir21         : out std_logic;
      iob21        : in  std_logic;
      i21          : in  std_logic;
      i20          : in  std_logic;
      iob20        : in  std_logic;
      ir20         : out std_logic;
      ir19         : out std_logic;
      iob19        : in  std_logic;
      i19          : in  std_logic;
      i18          : in  std_logic;
      iob18        : in  std_logic;
      ir18         : out std_logic;
      ir17         : out std_logic;
      iob17        : in  std_logic;
      i17          : in  std_logic;
      i16          : in  std_logic;
      iob16        : in  std_logic;
      ir16         : out std_logic;
      \-destimod1\ : in  std_logic;
      i48          : in  std_logic;
      ir48         : out std_logic;
      ir47         : out std_logic;
      iob47        : in  std_logic;
      i47          : in  std_logic;
      i46          : in  std_logic;
      iob46        : in  std_logic;
      ir46         : out std_logic;
      ir45         : out std_logic;
      iob45        : in  std_logic;
      i45          : in  std_logic;
      i44          : in  std_logic;
      iob44        : in  std_logic;
      ir44         : out std_logic;
      ir43         : out std_logic;
      iob43        : in  std_logic;
      i43          : in  std_logic;
      i42          : in  std_logic;
      iob42        : in  std_logic;
      ir42         : out std_logic;
      ir41         : out std_logic;
      iob41        : in  std_logic;
      i41          : in  std_logic;
      i40          : in  std_logic;
      iob40        : in  std_logic;
      ir40         : out std_logic;
      ir39         : out std_logic;
      iob39        : in  std_logic;
      i39          : in  std_logic;
      i38          : in  std_logic;
      iob38        : in  std_logic;
      ir38         : out std_logic;
      ir37         : out std_logic;
      iob37        : in  std_logic;
      i37          : in  std_logic;
      i36          : in  std_logic;
      iob36        : in  std_logic;
      ir36         : out std_logic;
      ir35         : out std_logic;
      iob35        : in  std_logic;
      i35          : in  std_logic;
      i34          : in  std_logic;
      iob34        : in  std_logic;
      ir34         : out std_logic;
      ir33         : out std_logic;
      iob33        : in  std_logic;
      i33          : in  std_logic;
      i32          : in  std_logic;
      iob32        : in  std_logic;
      ir32         : out std_logic;
      ir31         : out std_logic;
      iob31        : in  std_logic;
      i31          : in  std_logic;
      i30          : in  std_logic;
      iob30        : in  std_logic;
      ir30         : out std_logic;
      ir29         : out std_logic;
      iob29        : in  std_logic;
      i29          : in  std_logic;
      i28          : in  std_logic;
      iob28        : in  std_logic;
      ir28         : out std_logic;
      ir27         : out std_logic;
      iob27        : in  std_logic;
      i27          : in  std_logic;
      i26          : in  std_logic;
      iob26        : in  std_logic;
      ir26         : out std_logic;
      ir25         : out std_logic;
      iob25        : in  std_logic;
      i25          : in  std_logic;
      i24          : in  std_logic;
      iob24        : in  std_logic;
      ir24         : out std_logic
      );
  end component;

  component cadr_iwr is
    port (
      iwr47 : out std_logic;
      aa15  : in  std_logic;
      aa14  : in  std_logic;
      iwr46 : out std_logic;
      iwr45 : out std_logic;
      aa13  : in  std_logic;
      aa12  : in  std_logic;
      iwr44 : out std_logic;
      clk2c : in  std_logic;
      iwr43 : out std_logic;
      aa11  : in  std_logic;
      aa10  : in  std_logic;
      iwr42 : out std_logic;
      iwr41 : out std_logic;
      aa9   : in  std_logic;
      aa8   : in  std_logic;
      iwr40 : out std_logic;
      iwr39 : out std_logic;
      aa7   : in  std_logic;
      aa6   : in  std_logic;
      iwr38 : out std_logic;
      iwr37 : out std_logic;
      aa5   : in  std_logic;
      aa4   : in  std_logic;
      iwr36 : out std_logic;
      iwr35 : out std_logic;
      aa3   : in  std_logic;
      aa2   : in  std_logic;
      iwr34 : out std_logic;
      iwr33 : out std_logic;
      aa1   : in  std_logic;
      aa0   : in  std_logic;
      iwr32 : out std_logic;
      iwr15 : out std_logic;
      m15   : in  std_logic;
      m14   : in  std_logic;
      iwr14 : out std_logic;
      iwr13 : out std_logic;
      m13   : in  std_logic;
      m12   : in  std_logic;
      iwr12 : out std_logic;
      clk4c : in  std_logic;
      iwr11 : out std_logic;
      m11   : in  std_logic;
      m10   : in  std_logic;
      iwr10 : out std_logic;
      iwr9  : out std_logic;
      m9    : in  std_logic;
      m8    : in  std_logic;
      iwr8  : out std_logic;
      iwr7  : out std_logic;
      m7    : in  std_logic;
      m6    : in  std_logic;
      iwr6  : out std_logic;
      iwr5  : out std_logic;
      m5    : in  std_logic;
      m4    : in  std_logic;
      iwr4  : out std_logic;
      iwr3  : out std_logic;
      m3    : in  std_logic;
      m2    : in  std_logic;
      iwr2  : out std_logic;
      iwr1  : out std_logic;
      m1    : in  std_logic;
      m0    : in  std_logic;
      iwr0  : out std_logic;
      iwr31 : out std_logic;
      m31   : in  std_logic;
      m30   : in  std_logic;
      iwr30 : out std_logic;
      iwr29 : out std_logic;
      m29   : in  std_logic;
      m28   : in  std_logic;
      iwr28 : out std_logic;
      iwr27 : out std_logic;
      m27   : in  std_logic;
      m26   : in  std_logic;
      iwr26 : out std_logic;
      iwr25 : out std_logic;
      m25   : in  std_logic;
      m24   : in  std_logic;
      iwr24 : out std_logic;
      iwr23 : out std_logic;
      m23   : in  std_logic;
      m22   : in  std_logic;
      iwr22 : out std_logic;
      iwr21 : out std_logic;
      m21   : in  std_logic;
      m20   : in  std_logic;
      iwr20 : out std_logic;
      iwr19 : out std_logic;
      m19   : in  std_logic;
      m18   : in  std_logic;
      iwr18 : out std_logic;
      iwr17 : out std_logic;
      m17   : in  std_logic;
      m16   : in  std_logic;
      iwr16 : out std_logic
      );
  end component;

  component cadr_l is
    port (
      l7         : out std_logic;
      ob7        : in  std_logic;
      ob6        : in  std_logic;
      l6         : out std_logic;
      l5         : out std_logic;
      ob5        : in  std_logic;
      ob4        : in  std_logic;
      l4         : out std_logic;
      clk3f      : in  std_logic;
      l3         : out std_logic;
      ob3        : in  std_logic;
      ob2        : in  std_logic;
      l2         : out std_logic;
      l1         : out std_logic;
      ob1        : in  std_logic;
      ob0        : in  std_logic;
      l0         : out std_logic;
      l15        : out std_logic;
      ob15       : in  std_logic;
      ob14       : in  std_logic;
      l14        : out std_logic;
      l13        : out std_logic;
      ob13       : in  std_logic;
      ob12       : in  std_logic;
      l12        : out std_logic;
      l11        : out std_logic;
      ob11       : in  std_logic;
      ob10       : in  std_logic;
      l10        : out std_logic;
      l9         : out std_logic;
      ob9        : in  std_logic;
      ob8        : in  std_logic;
      l8         : out std_logic;
      l23        : out std_logic;
      ob23       : in  std_logic;
      ob22       : in  std_logic;
      l22        : out std_logic;
      l21        : out std_logic;
      ob21       : in  std_logic;
      ob20       : in  std_logic;
      l20        : out std_logic;
      l19        : out std_logic;
      ob19       : in  std_logic;
      ob18       : in  std_logic;
      l18        : out std_logic;
      l17        : out std_logic;
      ob17       : in  std_logic;
      ob16       : in  std_logic;
      l16        : out std_logic;
      l31        : out std_logic;
      ob31       : in  std_logic;
      ob30       : in  std_logic;
      l30        : out std_logic;
      l29        : out std_logic;
      ob29       : in  std_logic;
      ob28       : in  std_logic;
      l28        : out std_logic;
      l27        : out std_logic;
      ob27       : in  std_logic;
      ob26       : in  std_logic;
      l26        : out std_logic;
      l25        : out std_logic;
      ob25       : in  std_logic;
      ob24       : in  std_logic;
      lparl      : out std_logic;
      \-lparm\   : out std_logic;
      lparity    : out std_logic;
      \-lparity\ : out std_logic;
      l24        : out std_logic
      );
  end component;

  component cadr_lc is
    port (
      \-lcdrive\          : out std_logic;
      needfetch           : in  std_logic;
      mf24                : out std_logic;
      mf25                : out std_logic;
      \lc byte mode\      : in  std_logic;
      mf26                : out std_logic;
      \prog.unibus.reset\ : in  std_logic;
      mf27                : out std_logic;
      \int.enable\        : in  std_logic;
      mf28                : out std_logic;
      \sequence.break\    : in  std_logic;
      mf29                : out std_logic;
      lc25                : out std_logic;
      mf30                : out std_logic;
      lc24                : out std_logic;
      mf31                : out std_logic;
      lcdrive             : out std_logic;
      srclc               : out std_logic;
      tse1a               : in  std_logic;
      lc7                 : out std_logic;
      mf0                 : out std_logic;
      lc6                 : out std_logic;
      mf1                 : out std_logic;
      lc5                 : out std_logic;
      mf2                 : out std_logic;
      lc4                 : out std_logic;
      mf3                 : out std_logic;
      lc3                 : in  std_logic;
      mf4                 : out std_logic;
      lc2                 : in  std_logic;
      mf5                 : out std_logic;
      lc1                 : in  std_logic;
      mf6                 : out std_logic;
      lc0b                : in  std_logic;
      mf7                 : out std_logic;
      lc23                : out std_logic;
      mf16                : out std_logic;
      lc22                : out std_logic;
      mf17                : out std_logic;
      lc21                : out std_logic;
      mf18                : out std_logic;
      lc20                : out std_logic;
      mf19                : out std_logic;
      lc19                : out std_logic;
      mf20                : out std_logic;
      lc18                : out std_logic;
      mf21                : out std_logic;
      lc17                : out std_logic;
      mf22                : out std_logic;
      lc16                : out std_logic;
      mf23                : out std_logic;
      lc15                : out std_logic;
      mf8                 : out std_logic;
      lc14                : out std_logic;
      mf9                 : out std_logic;
      lc13                : out std_logic;
      mf10                : out std_logic;
      lc12                : out std_logic;
      mf11                : out std_logic;
      lc11                : out std_logic;
      mf12                : out std_logic;
      lc10                : out std_logic;
      mf13                : out std_logic;
      lc9                 : out std_logic;
      mf14                : out std_logic;
      lc8                 : out std_logic;
      mf15                : out std_logic;
      clk1a               : in  std_logic;
      ob20                : in  std_logic;
      ob21                : in  std_logic;
      ob22                : in  std_logic;
      ob23                : in  std_logic;
      \-destlc\           : in  std_logic;
      \-lcry19\           : out std_logic;
      \-lcry23\           : out std_logic;
      ob16                : in  std_logic;
      ob17                : in  std_logic;
      ob18                : in  std_logic;
      ob19                : in  std_logic;
      \-lcry15\           : out std_logic;
      clk2a               : in  std_logic;
      ob12                : in  std_logic;
      ob13                : in  std_logic;
      ob14                : in  std_logic;
      ob15                : in  std_logic;
      \-lcry11\           : out std_logic;
      clk2c               : in  std_logic;
      ob8                 : in  std_logic;
      ob9                 : in  std_logic;
      ob10                : in  std_logic;
      ob11                : in  std_logic;
      \-srclc\            : in  std_logic;
      ob24                : in  std_logic;
      ob25                : in  std_logic;
      ob4                 : in  std_logic;
      ob5                 : in  std_logic;
      ob6                 : in  std_logic;
      ob7                 : in  std_logic;
      \-lcry3\            : in  std_logic;
      \-lcry7\            : out std_logic
      );
  end component;

  component cadr_lcc is
    port (
      \lc byte mode\               : in  std_logic;
      \-lcinc\                     : out std_logic;
      lca1                         : out std_logic;
      lc1                          : out std_logic;
      lca0                         : out std_logic;
      lc0                          : out std_logic;
      lcinc                        : out std_logic;
      lcry3                        : out std_logic;
      lca3                         : out std_logic;
      lc3                          : out std_logic;
      lca2                         : out std_logic;
      lc2                          : out std_logic;
      \-destlc\                    : in  std_logic;
      ob3                          : in  std_logic;
      ob2                          : in  std_logic;
      clk2a                        : in  std_logic;
      ob1                          : in  std_logic;
      ob0                          : in  std_logic;
      lc0b                         : out std_logic;
      \inst in left half\          : out std_logic;
      \-ir4\                       : in  std_logic;
      \-sh4\                       : out std_logic;
      \-sh3\                       : out std_logic;
      \-ir3\                       : in  std_logic;
      \inst in 2nd or 4th quarter\ : out std_logic;
      \-lc modifies mrot\          : out std_logic;
      spc14                        : in  std_logic;
      \-srcspcpopreal\             : in  std_logic;
      \-ifetch\                    : out std_logic;
      needfetch                    : out std_logic;
      \have wrong word\            : out std_logic;
      \last byte in word\          : out std_logic;
      ir10                         : in  std_logic;
      ir11                         : in  std_logic;
      \-newlc\                     : out std_logic;
      \-newlc.in\                  : out std_logic;
      \-reset\                     : in  std_logic;
      newlc                        : out std_logic;
      int                          : in  std_logic;
      sintr                        : out std_logic;
      clk3c                        : in  std_logic;
      \next.instrd\                : out std_logic;
      \next.instr\                 : out std_logic;
      \-spop\                      : in  std_logic;
      \-needfetch\                 : out std_logic;
      spcmung                      : out std_logic;
      ir24                         : in  std_logic;
      irdisp                       : in  std_logic;
      spc1                         : in  std_logic;
      spc1a                        : out std_logic
      );
  end component;

  component cadr_lpc is
    port (
      pc8        : in  std_logic;
      pc9        : in  std_logic;
      pc10       : in  std_logic;
      pc13b      : out std_logic;
      pc11       : in  std_logic;
      pc12b      : out std_logic;
      pc12       : in  std_logic;
      pc11b      : out std_logic;
      pc13       : in  std_logic;
      pc10b      : out std_logic;
      pc9b       : out std_logic;
      pc8b       : out std_logic;
      pc0        : in  std_logic;
      pc7b       : out std_logic;
      pc1        : in  std_logic;
      pc6b       : out std_logic;
      pc2        : in  std_logic;
      pc5b       : out std_logic;
      pc3        : in  std_logic;
      pc4b       : out std_logic;
      pc4        : in  std_logic;
      pc3b       : out std_logic;
      pc5        : in  std_logic;
      pc2b       : out std_logic;
      pc6        : in  std_logic;
      pc1b       : out std_logic;
      pc7        : in  std_logic;
      pc0b       : out std_logic;
      irdisp     : in  std_logic;
      ir25       : in  std_logic;
      wpc12      : out std_logic;
      lpc13      : out std_logic;
      wpc13      : out std_logic;
      lpc8       : out std_logic;
      wpc8       : out std_logic;
      lpc9       : out std_logic;
      wpc9       : out std_logic;
      wpc10      : out std_logic;
      lpc10      : out std_logic;
      wpc11      : out std_logic;
      lpc11      : out std_logic;
      lpc4       : out std_logic;
      wpc4       : out std_logic;
      lpc5       : out std_logic;
      wpc5       : out std_logic;
      wpc6       : out std_logic;
      lpc6       : out std_logic;
      wpc7       : out std_logic;
      lpc7       : out std_logic;
      lpc0       : out std_logic;
      wpc0       : out std_logic;
      lpc1       : out std_logic;
      wpc1       : out std_logic;
      wpc2       : out std_logic;
      lpc2       : out std_logic;
      wpc3       : out std_logic;
      lpc3       : out std_logic;
      \lpc.hold\ : in  std_logic;
      clk4b      : in  std_logic;
      lpc12      : out std_logic
      );
  end component;

  component cadr_mctl is
    port (
      clk4e      : in  std_logic;
      wadr4      : in  std_logic;
      ir30       : in  std_logic;
      \-madr4a\  : out std_logic;
      \-madr4b\  : out std_logic;
      wadr0      : in  std_logic;
      ir26       : in  std_logic;
      \-madr0b\  : out std_logic;
      wadr1      : in  std_logic;
      ir27       : in  std_logic;
      \-madr1b\  : out std_logic;
      \-madr2b\  : out std_logic;
      ir28       : in  std_logic;
      wadr2      : in  std_logic;
      \-madr3b\  : out std_logic;
      ir29       : in  std_logic;
      wadr3      : in  std_logic;
      mmem15     : out std_logic;
      mmem14     : out std_logic;
      mmem13     : out std_logic;
      mmem12     : out std_logic;
      mmem11     : out std_logic;
      mmem10     : out std_logic;
      mmem9      : out std_logic;
      mmem8      : out std_logic;
      mmem7      : out std_logic;
      mmem6      : out std_logic;
      mmem5      : out std_logic;
      mmem4      : out std_logic;
      mmem3      : out std_logic;
      mmem2      : out std_logic;
      mmem1      : out std_logic;
      mmem0      : out std_logic;
      mpass      : out std_logic;
      tse4a      : in  std_logic;
      srcm       : out std_logic;
      \-ir31\    : in  std_logic;
      \-mpass\   : out std_logic;
      mpassl     : out std_logic;
      \-mpassm\  : out std_logic;
      \-mpassl\  : out std_logic;
      destmd     : in  std_logic;
      \-madr0a\  : out std_logic;
      \-madr1a\  : out std_logic;
      \-madr2a\  : out std_logic;
      \-madr3a\  : out std_logic;
      mmemparity : out std_logic;
      mmem31     : out std_logic;
      mmem30     : out std_logic;
      mmem29     : out std_logic;
      mmem28     : out std_logic;
      mmem27     : out std_logic;
      mmem26     : out std_logic;
      mmem25     : out std_logic;
      mmem24     : out std_logic;
      mmem23     : out std_logic;
      mmem22     : out std_logic;
      mmem21     : out std_logic;
      mmem20     : out std_logic;
      mmem19     : out std_logic;
      mmem18     : out std_logic;
      mmem17     : out std_logic;
      mmem16     : out std_logic;
      wp4b       : in  std_logic;
      \-mwpa\    : out std_logic;
      \-mwpb\    : out std_logic
      );
  end component;

  component cadr_md is
    port (
      \-mddrive\  : out std_logic;
      \-md31\     : out std_logic;
      mf24        : out std_logic;
      \-md30\     : out std_logic;
      mf25        : out std_logic;
      \-md29\     : out std_logic;
      mf26        : out std_logic;
      \-md28\     : out std_logic;
      mf27        : out std_logic;
      \-md27\     : out std_logic;
      mf28        : out std_logic;
      \-md26\     : out std_logic;
      mf29        : out std_logic;
      \-md25\     : out std_logic;
      mf30        : out std_logic;
      \-md24\     : out std_logic;
      mf31        : out std_logic;
      \-md23\     : out std_logic;
      mf16        : out std_logic;
      \-md22\     : out std_logic;
      mf17        : out std_logic;
      \-md21\     : out std_logic;
      mf18        : out std_logic;
      \-md20\     : out std_logic;
      mf19        : out std_logic;
      \-md19\     : out std_logic;
      mf20        : out std_logic;
      \-md18\     : out std_logic;
      mf21        : out std_logic;
      \-md17\     : out std_logic;
      mf22        : out std_logic;
      \-md16\     : out std_logic;
      mf23        : out std_logic;
      \-md7\      : out std_logic;
      mf0         : out std_logic;
      \-md6\      : out std_logic;
      mf1         : out std_logic;
      \-md5\      : out std_logic;
      mf2         : out std_logic;
      \-md4\      : out std_logic;
      mf3         : out std_logic;
      \-md3\      : out std_logic;
      mf4         : out std_logic;
      \-md2\      : out std_logic;
      mf5         : out std_logic;
      \-md1\      : out std_logic;
      mf6         : out std_logic;
      \-md0\      : out std_logic;
      mf7         : out std_logic;
      srcmd       : out std_logic;
      tse2        : in  std_logic;
      \-md15\     : out std_logic;
      mf8         : out std_logic;
      \-md14\     : out std_logic;
      mf9         : out std_logic;
      \-md13\     : out std_logic;
      mf10        : out std_logic;
      \-md12\     : out std_logic;
      mf11        : out std_logic;
      \-md11\     : out std_logic;
      mf12        : out std_logic;
      \-md10\     : out std_logic;
      mf13        : out std_logic;
      \-md9\      : out std_logic;
      mf14        : out std_logic;
      \-md8\      : out std_logic;
      mf15        : out std_logic;
      \-mds31\    : in  std_logic;
      \-mds30\    : in  std_logic;
      \-mds29\    : in  std_logic;
      \-mds28\    : in  std_logic;
      mdclk       : out std_logic;
      \-mds27\    : in  std_logic;
      \-mds26\    : in  std_logic;
      \-mds25\    : in  std_logic;
      \-mds24\    : in  std_logic;
      \-mds7\     : in  std_logic;
      \-mds6\     : in  std_logic;
      \-mds5\     : in  std_logic;
      \-mds4\     : in  std_logic;
      \-mds3\     : in  std_logic;
      \-mds2\     : in  std_logic;
      \-mds1\     : in  std_logic;
      \-mds0\     : in  std_logic;
      \-mds23\    : in  std_logic;
      \-mds22\    : in  std_logic;
      \-mds21\    : in  std_logic;
      \-mds20\    : in  std_logic;
      \-mds19\    : in  std_logic;
      \-mds18\    : in  std_logic;
      \-mds17\    : in  std_logic;
      \-mds16\    : in  std_logic;
      destmdr     : out std_logic;
      \-clk2c\    : in  std_logic;
      loadmd      : out std_logic;
      \-loadmd\   : in  std_logic;
      \-destmdr\  : in  std_logic;
      \-mds15\    : in  std_logic;
      \-mds14\    : in  std_logic;
      \-mds13\    : in  std_logic;
      \-mds12\    : in  std_logic;
      \-mds11\    : in  std_logic;
      \-mds10\    : in  std_logic;
      \-mds9\     : in  std_logic;
      \-mds8\     : in  std_logic;
      mdgetspar   : out std_logic;
      \-ignpar\   : in  std_logic;
      mdhaspar    : out std_logic;
      \mempar in\ : in  std_logic;
      mdpar       : out std_logic;
      \-srcmd\    : in  std_logic
      );
  end component;

  component cadr_mds is
    port (
      \-memdrive.a\ : in  std_logic;
      \-md31\       : in  std_logic;
      mem24         : out std_logic;
      \-md30\       : in  std_logic;
      mem25         : out std_logic;
      \-md29\       : in  std_logic;
      mem26         : out std_logic;
      \-md28\       : in  std_logic;
      \-md27\       : in  std_logic;
      mem28         : out std_logic;
      \-md26\       : in  std_logic;
      mem29         : out std_logic;
      \-md25\       : in  std_logic;
      mem30         : out std_logic;
      \-md24\       : in  std_logic;
      mem31         : out std_logic;
      \-memdrive.b\ : in  std_logic;
      \-md7\        : in  std_logic;
      mem0          : out std_logic;
      \-md6\        : in  std_logic;
      mem1          : out std_logic;
      \-md5\        : in  std_logic;
      mem2          : out std_logic;
      \-md4\        : in  std_logic;
      mem3          : out std_logic;
      \-md3\        : in  std_logic;
      mem4          : out std_logic;
      \-md2\        : in  std_logic;
      mem5          : out std_logic;
      \-md1\        : in  std_logic;
      mem6          : out std_logic;
      \-md0\        : in  std_logic;
      mem7          : out std_logic;
      \-md23\       : in  std_logic;
      mem16         : out std_logic;
      \-md22\       : in  std_logic;
      mem17         : out std_logic;
      \-md21\       : in  std_logic;
      mem18         : out std_logic;
      \-md20\       : in  std_logic;
      mem19         : out std_logic;
      \-md19\       : in  std_logic;
      mem20         : out std_logic;
      \-md18\       : in  std_logic;
      mem21         : out std_logic;
      \-md17\       : in  std_logic;
      mem22         : out std_logic;
      \-md16\       : in  std_logic;
      mem23         : out std_logic;
      \-md15\       : in  std_logic;
      mem8          : out std_logic;
      \-md14\       : in  std_logic;
      mem9          : out std_logic;
      \-md13\       : in  std_logic;
      mem10         : out std_logic;
      \-md12\       : in  std_logic;
      mem11         : out std_logic;
      \-md11\       : in  std_logic;
      mem12         : out std_logic;
      \-md10\       : in  std_logic;
      mem13         : out std_logic;
      \-md9\        : in  std_logic;
      mem14         : out std_logic;
      \-md8\        : in  std_logic;
      mem15         : out std_logic;
      mdsela        : in  std_logic;
      ob20          : in  std_logic;
      \-mds20\      : out std_logic;
      ob21          : in  std_logic;
      \-mds21\      : out std_logic;
      \-mds22\      : out std_logic;
      ob22          : in  std_logic;
      \-mds23\      : out std_logic;
      ob23          : in  std_logic;
      ob28          : in  std_logic;
      \-mds28\      : out std_logic;
      ob29          : in  std_logic;
      \-mds29\      : out std_logic;
      \-mds30\      : out std_logic;
      ob30          : in  std_logic;
      \-mds31\      : out std_logic;
      ob31          : in  std_logic;
      mdparodd      : in  std_logic;
      \mempar out\  : out std_logic;
      mdselb        : in  std_logic;
      ob12          : in  std_logic;
      \-mds12\      : out std_logic;
      ob13          : in  std_logic;
      \-mds13\      : out std_logic;
      \-mds14\      : out std_logic;
      ob14          : in  std_logic;
      \-mds15\      : out std_logic;
      ob15          : in  std_logic;
      ob16          : in  std_logic;
      \-mds16\      : out std_logic;
      ob17          : in  std_logic;
      \-mds17\      : out std_logic;
      \-mds18\      : out std_logic;
      ob18          : in  std_logic;
      \-mds19\      : out std_logic;
      ob19          : in  std_logic;
      ob8           : in  std_logic;
      \-mds8\       : out std_logic;
      ob9           : in  std_logic;
      \-mds9\       : out std_logic;
      \-mds10\      : out std_logic;
      ob10          : in  std_logic;
      \-mds11\      : out std_logic;
      ob11          : in  std_logic;
      ob0           : in  std_logic;
      \-mds0\       : out std_logic;
      ob1           : in  std_logic;
      \-mds1\       : out std_logic;
      \-mds2\       : out std_logic;
      ob2           : in  std_logic;
      \-mds3\       : out std_logic;
      ob3           : in  std_logic;
      ob4           : in  std_logic;
      \-mds4\       : out std_logic;
      ob5           : in  std_logic;
      \-mds5\       : out std_logic;
      \-mds6\       : out std_logic;
      ob6           : in  std_logic;
      \-mds7\       : out std_logic;
      ob7           : in  std_logic;
      ob24          : in  std_logic;
      \-mds24\      : out std_logic;
      ob25          : in  std_logic;
      \-mds25\      : out std_logic;
      \-mds26\      : out std_logic;
      ob26          : in  std_logic;
      \-mds27\      : out std_logic;
      ob27          : in  std_logic;
      mem27         : out std_logic
      );
  end component;

  component cadr_mf is
    port (
      tse1a      : in  std_logic;
      mfenb      : out std_logic;
      \-mfdrive\ : out std_logic;
      mf23       : in  std_logic;
      m16        : out std_logic;
      mf22       : in  std_logic;
      m17        : out std_logic;
      mf21       : in  std_logic;
      m18        : out std_logic;
      mf20       : in  std_logic;
      m19        : out std_logic;
      mf19       : in  std_logic;
      m20        : out std_logic;
      mf18       : in  std_logic;
      m21        : out std_logic;
      mf17       : in  std_logic;
      m22        : out std_logic;
      mf16       : in  std_logic;
      m23        : out std_logic;
      mfdrive    : out std_logic;
      mf15       : in  std_logic;
      m8         : out std_logic;
      mf14       : in  std_logic;
      m9         : out std_logic;
      mf13       : in  std_logic;
      m10        : out std_logic;
      mf12       : in  std_logic;
      m11        : out std_logic;
      mf11       : in  std_logic;
      m12        : out std_logic;
      mf10       : in  std_logic;
      m13        : out std_logic;
      mf9        : in  std_logic;
      m14        : out std_logic;
      mf8        : in  std_logic;
      m15        : out std_logic;
      mf7        : in  std_logic;
      m0         : out std_logic;
      mf6        : in  std_logic;
      m1         : out std_logic;
      mf5        : in  std_logic;
      m2         : out std_logic;
      mf4        : in  std_logic;
      m3         : out std_logic;
      mf3        : in  std_logic;
      m4         : out std_logic;
      mf2        : in  std_logic;
      m5         : out std_logic;
      mf1        : in  std_logic;
      m6         : out std_logic;
      mf0        : in  std_logic;
      m7         : out std_logic;
      mf31       : in  std_logic;
      m24        : out std_logic;
      mf30       : in  std_logic;
      m25        : out std_logic;
      mf29       : in  std_logic;
      m26        : out std_logic;
      mf28       : in  std_logic;
      m27        : out std_logic;
      mf27       : in  std_logic;
      m28        : out std_logic;
      mf26       : in  std_logic;
      m29        : out std_logic;
      mf25       : in  std_logic;
      m30        : out std_logic;
      mf24       : in  std_logic;
      m31        : out std_logic;
      pdlenb     : in  std_logic;
      spcenb     : in  std_logic;
      \-srcm\    : out std_logic;
      \-ir31\    : in  std_logic;
      \-mpass\   : in  std_logic
      );
  end component;

  component cadr_mlatch is
    port (
      \-mpassm\  : in  std_logic;
      m23        : out std_logic;
      mmem23     : in  std_logic;
      mmem22     : out std_logic;
      m22        : out std_logic;
      m21        : out std_logic;
      mmem21     : in  std_logic;
      mmem20     : out std_logic;
      m20        : out std_logic;
      clk4a      : in  std_logic;
      m19        : out std_logic;
      mmem19     : in  std_logic;
      mmem18     : out std_logic;
      m18        : out std_logic;
      m17        : out std_logic;
      mmem17     : in  std_logic;
      mmem16     : out std_logic;
      m16        : out std_logic;
      m15        : out std_logic;
      mmem15     : in  std_logic;
      mmem14     : out std_logic;
      m14        : out std_logic;
      m13        : out std_logic;
      mmem13     : in  std_logic;
      mmem12     : out std_logic;
      m12        : out std_logic;
      m11        : out std_logic;
      mmem11     : in  std_logic;
      mmem10     : out std_logic;
      m10        : out std_logic;
      m9         : out std_logic;
      mmem9      : in  std_logic;
      mmem8      : out std_logic;
      m8         : out std_logic;
      m7         : out std_logic;
      mmem7      : in  std_logic;
      mmem6      : out std_logic;
      m6         : out std_logic;
      m5         : out std_logic;
      mmem5      : in  std_logic;
      mmem4      : out std_logic;
      m4         : out std_logic;
      m3         : out std_logic;
      mmem3      : in  std_logic;
      mmem2      : in  std_logic;
      m2         : out std_logic;
      m1         : out std_logic;
      mmem1      : out std_logic;
      mmem0      : out std_logic;
      m0         : out std_logic;
      \-mpassl\  : in  std_logic;
      l15        : in  std_logic;
      mf8        : out std_logic;
      l14        : in  std_logic;
      mf9        : out std_logic;
      l13        : in  std_logic;
      mf10       : out std_logic;
      l12        : in  std_logic;
      mf11       : out std_logic;
      l11        : in  std_logic;
      mf12       : out std_logic;
      l10        : in  std_logic;
      mf13       : out std_logic;
      l9         : in  std_logic;
      mf14       : out std_logic;
      l8         : in  std_logic;
      mf15       : out std_logic;
      mpassl     : in  std_logic;
      l7         : in  std_logic;
      mf0        : out std_logic;
      l6         : in  std_logic;
      mf1        : out std_logic;
      l5         : in  std_logic;
      mf2        : out std_logic;
      l4         : in  std_logic;
      mf3        : out std_logic;
      l3         : in  std_logic;
      mf4        : out std_logic;
      l2         : in  std_logic;
      mf5        : out std_logic;
      l1         : in  std_logic;
      mf6        : out std_logic;
      l0         : in  std_logic;
      mf7        : out std_logic;
      mmemparity : out std_logic;
      mparity    : out std_logic;
      m31        : out std_logic;
      mmem31     : in  std_logic;
      mmem30     : out std_logic;
      m30        : out std_logic;
      m29        : out std_logic;
      mmem29     : in  std_logic;
      mmem28     : out std_logic;
      m28        : out std_logic;
      m27        : out std_logic;
      mmem27     : in  std_logic;
      mmem26     : out std_logic;
      m26        : out std_logic;
      m25        : out std_logic;
      mmem25     : in  std_logic;
      mmem24     : out std_logic;
      m24        : out std_logic;
      l31        : in  std_logic;
      mf24       : out std_logic;
      l30        : in  std_logic;
      mf25       : out std_logic;
      l29        : in  std_logic;
      mf26       : out std_logic;
      l28        : in  std_logic;
      mf27       : out std_logic;
      l27        : in  std_logic;
      mf28       : out std_logic;
      l26        : in  std_logic;
      mf29       : out std_logic;
      l25        : in  std_logic;
      mf30       : out std_logic;
      l24        : in  std_logic;
      mf31       : out std_logic;
      l23        : in  std_logic;
      mf16       : out std_logic;
      l22        : in  std_logic;
      mf17       : out std_logic;
      l21        : in  std_logic;
      mf18       : out std_logic;
      l20        : in  std_logic;
      mf19       : out std_logic;
      l19        : in  std_logic;
      mf20       : out std_logic;
      l18        : in  std_logic;
      mf21       : out std_logic;
      l17        : in  std_logic;
      mf22       : out std_logic;
      l16        : in  std_logic;
      mf23       : out std_logic
      );
  end component;

  component cadr_mmem is
    port (
      \-mwpa\    : in  std_logic;
      l16        : in  std_logic;
      \-madr4a\  : in  std_logic;
      mmem16     : out std_logic;
      mmem17     : out std_logic;
      \-madr3a\  : in  std_logic;
      \-madr2a\  : in  std_logic;
      \-madr1a\  : in  std_logic;
      \-madr0a\  : in  std_logic;
      l17        : in  std_logic;
      \-mwpb\    : in  std_logic;
      l12        : in  std_logic;
      \-madr4b\  : in  std_logic;
      mmem12     : out std_logic;
      mmem13     : out std_logic;
      \-madr3b\  : in  std_logic;
      \-madr2b\  : in  std_logic;
      \-madr1b\  : in  std_logic;
      \-madr0b\  : in  std_logic;
      l13        : in  std_logic;
      l8         : in  std_logic;
      mmem8      : out std_logic;
      mmem9      : out std_logic;
      l9         : in  std_logic;
      l4         : in  std_logic;
      mmem4      : out std_logic;
      mmem5      : out std_logic;
      l5         : in  std_logic;
      l0         : in  std_logic;
      mmem0      : out std_logic;
      mmem1      : out std_logic;
      l1         : in  std_logic;
      l18        : in  std_logic;
      mmem18     : out std_logic;
      mmem19     : out std_logic;
      l19        : in  std_logic;
      l14        : in  std_logic;
      mmem14     : out std_logic;
      mmem15     : out std_logic;
      l15        : in  std_logic;
      l10        : in  std_logic;
      mmem10     : out std_logic;
      mmem11     : out std_logic;
      l11        : in  std_logic;
      l6         : in  std_logic;
      mmem6      : out std_logic;
      mmem7      : out std_logic;
      l7         : in  std_logic;
      l2         : in  std_logic;
      mmem2      : out std_logic;
      mmem3      : out std_logic;
      l3         : in  std_logic;
      l28        : in  std_logic;
      mmem28     : out std_logic;
      mmem29     : out std_logic;
      l29        : in  std_logic;
      l24        : in  std_logic;
      mmem24     : out std_logic;
      mmem25     : out std_logic;
      l25        : in  std_logic;
      l20        : in  std_logic;
      mmem20     : out std_logic;
      mmem21     : out std_logic;
      l21        : in  std_logic;
      lparity    : in  std_logic;
      mmemparity : out std_logic;
      l30        : in  std_logic;
      mmem30     : out std_logic;
      mmem31     : out std_logic;
      l31        : in  std_logic;
      l26        : in  std_logic;
      mmem26     : out std_logic;
      mmem27     : out std_logic;
      l27        : in  std_logic;
      l22        : in  std_logic;
      mmem22     : out std_logic;
      mmem23     : out std_logic;
      l23        : in  std_logic
      );
  end component;

  component cadr_mo0 is
    port (
      alu15  : in  std_logic;
      r15    : in  std_logic;
      a15    : in  std_logic;
      ob15   : out std_logic;
      osel1b : in  std_logic;
      osel0b : in  std_logic;
      msk15  : in  std_logic;
      alu14  : in  std_logic;
      alu16  : in  std_logic;
      r14    : in  std_logic;
      a14    : in  std_logic;
      ob14   : out std_logic;
      msk14  : in  std_logic;
      alu13  : in  std_logic;
      r13    : in  std_logic;
      a13    : in  std_logic;
      ob13   : out std_logic;
      msk13  : in  std_logic;
      alu12  : in  std_logic;
      r12    : in  std_logic;
      a12    : in  std_logic;
      ob12   : out std_logic;
      msk12  : in  std_logic;
      alu11  : in  std_logic;
      alu7   : in  std_logic;
      r7     : in  std_logic;
      a7     : in  std_logic;
      ob7    : out std_logic;
      msk7   : in  std_logic;
      alu6   : in  std_logic;
      alu8   : in  std_logic;
      r6     : in  std_logic;
      a6     : in  std_logic;
      ob6    : out std_logic;
      msk6   : in  std_logic;
      alu5   : in  std_logic;
      r5     : in  std_logic;
      a5     : in  std_logic;
      ob5    : out std_logic;
      msk5   : in  std_logic;
      alu4   : in  std_logic;
      r4     : in  std_logic;
      a4     : in  std_logic;
      ob4    : out std_logic;
      msk4   : in  std_logic;
      alu3   : in  std_logic;
      r11    : in  std_logic;
      a11    : in  std_logic;
      ob11   : out std_logic;
      msk11  : in  std_logic;
      alu10  : in  std_logic;
      r10    : in  std_logic;
      a10    : in  std_logic;
      ob10   : out std_logic;
      msk10  : in  std_logic;
      alu9   : in  std_logic;
      r3     : in  std_logic;
      a3     : in  std_logic;
      ob3    : out std_logic;
      msk3   : in  std_logic;
      alu2   : in  std_logic;
      r2     : in  std_logic;
      a2     : in  std_logic;
      ob2    : out std_logic;
      msk2   : in  std_logic;
      r9     : in  std_logic;
      a9     : in  std_logic;
      ob9    : out std_logic;
      msk9   : in  std_logic;
      r8     : in  std_logic;
      a8     : in  std_logic;
      ob8    : out std_logic;
      msk8   : in  std_logic;
      r1     : in  std_logic;
      a1     : in  std_logic;
      ob1    : out std_logic;
      msk1   : in  std_logic;
      alu0   : in  std_logic;
      r0     : in  std_logic;
      a0     : in  std_logic;
      ob0    : out std_logic;
      msk0   : in  std_logic;
      q31    : in  std_logic;
      alu1   : in  std_logic
      );
  end component;

  component cadr_mo1 is
    port (
      alu31  : in  std_logic;
      r31    : in  std_logic;
      a31b   : in  std_logic;
      ob31   : out std_logic;
      osel1a : in  std_logic;
      osel0a : in  std_logic;
      msk31  : in  std_logic;
      alu30  : in  std_logic;
      alu32  : in  std_logic;
      r30    : in  std_logic;
      a30    : in  std_logic;
      ob30   : out std_logic;
      msk30  : in  std_logic;
      alu29  : in  std_logic;
      r29    : in  std_logic;
      a29    : in  std_logic;
      ob29   : out std_logic;
      msk29  : in  std_logic;
      alu28  : in  std_logic;
      r28    : in  std_logic;
      a28    : in  std_logic;
      ob28   : out std_logic;
      msk28  : in  std_logic;
      alu27  : in  std_logic;
      alu23  : in  std_logic;
      r23    : in  std_logic;
      a23    : in  std_logic;
      ob23   : out std_logic;
      msk23  : in  std_logic;
      alu22  : in  std_logic;
      alu24  : in  std_logic;
      r22    : in  std_logic;
      a22    : in  std_logic;
      ob22   : out std_logic;
      msk22  : in  std_logic;
      alu21  : in  std_logic;
      r21    : in  std_logic;
      a21    : in  std_logic;
      ob21   : out std_logic;
      msk21  : in  std_logic;
      alu20  : in  std_logic;
      r20    : in  std_logic;
      a20    : in  std_logic;
      ob20   : out std_logic;
      msk20  : in  std_logic;
      alu19  : in  std_logic;
      r27    : in  std_logic;
      a27    : in  std_logic;
      ob27   : out std_logic;
      msk27  : in  std_logic;
      alu26  : in  std_logic;
      r24    : in  std_logic;
      a24    : in  std_logic;
      ob24   : out std_logic;
      msk24  : in  std_logic;
      alu25  : in  std_logic;
      r26    : in  std_logic;
      a26    : in  std_logic;
      ob26   : out std_logic;
      msk26  : in  std_logic;
      r25    : in  std_logic;
      a25    : in  std_logic;
      ob25   : out std_logic;
      msk25  : in  std_logic;
      r19    : in  std_logic;
      a19    : in  std_logic;
      ob19   : out std_logic;
      msk19  : in  std_logic;
      alu18  : in  std_logic;
      r18    : in  std_logic;
      a18    : in  std_logic;
      ob18   : out std_logic;
      msk18  : in  std_logic;
      r17    : in  std_logic;
      a17    : in  std_logic;
      ob17   : out std_logic;
      msk17  : in  std_logic;
      alu16  : in  std_logic;
      r16    : in  std_logic;
      a16    : in  std_logic;
      ob16   : out std_logic;
      msk16  : in  std_logic;
      alu15  : in  std_logic;
      alu17  : in  std_logic
      );
  end component;

  component cadr_mskg4 is
    port (
      msk24   : out std_logic;
      msk25   : out std_logic;
      msk26   : out std_logic;
      msk27   : out std_logic;
      msk28   : out std_logic;
      msk29   : out std_logic;
      msk30   : out std_logic;
      msk31   : out std_logic;
      mskl0   : in  std_logic;
      mskl1   : in  std_logic;
      mskl2   : in  std_logic;
      mskl3   : in  std_logic;
      mskl4   : in  std_logic;
      mskr0   : in  std_logic;
      mskr1   : in  std_logic;
      mskr2   : in  std_logic;
      mskr3   : in  std_logic;
      mskr4   : in  std_logic;
      msk8    : out std_logic;
      msk9    : out std_logic;
      msk10   : out std_logic;
      msk11   : out std_logic;
      msk12   : out std_logic;
      msk13   : out std_logic;
      msk14   : out std_logic;
      msk15   : out std_logic;
      ir31    : in  std_logic;
      \-ir31\ : out std_logic;
      ir13    : in  std_logic;
      \-ir13\ : out std_logic;
      \-ir12\ : out std_logic;
      ir12    : in  std_logic;
      msk16   : out std_logic;
      msk17   : out std_logic;
      msk18   : out std_logic;
      msk19   : out std_logic;
      msk20   : out std_logic;
      msk21   : out std_logic;
      msk22   : out std_logic;
      msk23   : out std_logic;
      \a=m\   : out std_logic;
      msk1    : out std_logic;
      msk2    : out std_logic;
      msk3    : out std_logic;
      msk4    : out std_logic;
      msk5    : out std_logic;
      msk6    : out std_logic;
      msk7    : out std_logic;
      msk0    : out std_logic
      );
  end component;

  component cadr_npc is
    port (
      ipc13   : out std_logic;
      pc13    : out std_logic;
      ipc12   : out std_logic;
      pc12    : out std_logic;
      pccry11 : out std_logic;
      ipc9    : out std_logic;
      pc9     : out std_logic;
      ipc8    : out std_logic;
      pc8     : out std_logic;
      pccry7  : out std_logic;
      ipc11   : out std_logic;
      pc11    : out std_logic;
      ipc10   : out std_logic;
      pc10    : out std_logic;
      ipc5    : out std_logic;
      pc5     : out std_logic;
      pc4     : out std_logic;
      pccry3  : out std_logic;
      ipc7    : out std_logic;
      pc7     : out std_logic;
      ipc6    : out std_logic;
      pc6     : out std_logic;
      ipc1    : out std_logic;
      pc1     : out std_logic;
      ipc0    : out std_logic;
      pc0     : out std_logic;
      ipc3    : out std_logic;
      pc3     : out std_logic;
      ipc2    : out std_logic;
      pc2     : out std_logic;
      trapb   : in  std_logic;
      pcs1    : in  std_logic;
      dpc3    : out std_logic;
      ir15    : in  std_logic;
      spc3    : out std_logic;
      npc3    : out std_logic;
      npc2    : out std_logic;
      spc2    : out std_logic;
      ir14    : in  std_logic;
      dpc2    : out std_logic;
      pcs0    : in  std_logic;
      dpc1    : out std_logic;
      ir13    : in  std_logic;
      spc1a   : in  std_logic;
      npc1    : out std_logic;
      npc0    : out std_logic;
      spc0    : out std_logic;
      ir12    : in  std_logic;
      dpc0    : out std_logic;
      npc13   : out std_logic;
      npc12   : out std_logic;
      clk4b   : in  std_logic;
      npc11   : out std_logic;
      npc10   : out std_logic;
      npc9    : out std_logic;
      npc8    : out std_logic;
      npc7    : out std_logic;
      npc6    : out std_logic;
      npc5    : out std_logic;
      npc4    : out std_logic;
      trapa   : in  std_logic;
      dpc13   : out std_logic;
      ir25    : in  std_logic;
      spc13   : out std_logic;
      spc12   : out std_logic;
      ir24    : in  std_logic;
      dpc12   : out std_logic;
      dpc11   : out std_logic;
      ir23    : in  std_logic;
      spc11   : out std_logic;
      spc10   : out std_logic;
      ir22    : in  std_logic;
      dpc10   : out std_logic;
      dpc9    : out std_logic;
      ir21    : in  std_logic;
      spc9    : out std_logic;
      spc8    : out std_logic;
      ir20    : in  std_logic;
      dpc8    : out std_logic;
      dpc7    : out std_logic;
      ir19    : in  std_logic;
      spc7    : out std_logic;
      spc6    : out std_logic;
      ir18    : in  std_logic;
      dpc6    : out std_logic;
      dpc5    : out std_logic;
      ir17    : in  std_logic;
      spc5    : out std_logic;
      spc4    : out std_logic;
      ir16    : in  std_logic;
      dpc4    : in  std_logic;
      ipc4    : out std_logic
      );
  end component;

  component cadr_opcd is
    port (
      \-srcopc\       : in  std_logic;
      \-opcdrive\     : out std_logic;
      opc7            : in  std_logic;
      mf4             : out std_logic;
      opc6            : in  std_logic;
      mf5             : out std_logic;
      opc5            : in  std_logic;
      mf6             : out std_logic;
      opc4            : in  std_logic;
      mf7             : out std_logic;
      dc7             : in  std_logic;
      dc6             : in  std_logic;
      dc5             : in  std_logic;
      dc4             : in  std_logic;
      dcdrive         : out std_logic;
      opc3            : in  std_logic;
      mf0             : out std_logic;
      opc2            : in  std_logic;
      mf1             : out std_logic;
      opc1            : in  std_logic;
      mf2             : out std_logic;
      opc0            : in  std_logic;
      mf3             : out std_logic;
      dc3             : in  std_logic;
      dc2             : in  std_logic;
      dc1             : in  std_logic;
      dc0             : in  std_logic;
      tse1b           : in  std_logic;
      \-zero16.drive\ : out std_logic;
      zero16          : out std_logic;
      \zero16.drive\  : out std_logic;
      \zero12.drive\  : out std_logic;
      mf24            : out std_logic;
      mf25            : out std_logic;
      mf26            : out std_logic;
      mf27            : out std_logic;
      mf28            : out std_logic;
      mf29            : out std_logic;
      mf30            : out std_logic;
      mf31            : out std_logic;
      mf16            : out std_logic;
      mf17            : out std_logic;
      mf18            : out std_logic;
      mf19            : out std_logic;
      mf20            : out std_logic;
      mf21            : out std_logic;
      mf22            : out std_logic;
      mf23            : out std_logic;
      mf12            : out std_logic;
      mf13            : out std_logic;
      opc13           : in  std_logic;
      mf14            : out std_logic;
      opc12           : in  std_logic;
      mf15            : out std_logic;
      opc11           : in  std_logic;
      mf8             : out std_logic;
      opc10           : in  std_logic;
      mf9             : out std_logic;
      opc9            : in  std_logic;
      mf10            : out std_logic;
      opc8            : in  std_logic;
      mf11            : out std_logic;
      dc9             : in  std_logic;
      dc8             : in  std_logic;
      \-srcpdlidx\    : in  std_logic;
      \-srcpdlptr\    : in  std_logic;
      \-srcdc\        : in  std_logic
      );
  end component;

  component cadr_pdl0 is
    port (
      \-pdla0b\ : in  std_logic;
      \-pdla1b\ : in  std_logic;
      \-pdla2b\ : in  std_logic;
      \-pdla3b\ : in  std_logic;
      \-pdla4b\ : in  std_logic;
      pdlparity : out std_logic;
      \-pdla5b\ : in  std_logic;
      \-pdla6b\ : in  std_logic;
      \-pdla7b\ : in  std_logic;
      \-pdla8b\ : in  std_logic;
      \-pdla9b\ : in  std_logic;
      \-pwpa\   : in  std_logic;
      lparity   : in  std_logic;
      pdl28     : out std_logic;
      l28       : in  std_logic;
      pdl27     : out std_logic;
      l27       : in  std_logic;
      pdl26     : out std_logic;
      l26       : in  std_logic;
      pdl21     : out std_logic;
      \-pwpb\   : in  std_logic;
      l21       : in  std_logic;
      pdl20     : out std_logic;
      l20       : in  std_logic;
      pdl19     : out std_logic;
      l19       : in  std_logic;
      pdl18     : out std_logic;
      l18       : in  std_logic;
      pdl31     : out std_logic;
      l31       : in  std_logic;
      pdl30     : out std_logic;
      l30       : in  std_logic;
      pdl29     : out std_logic;
      l29       : in  std_logic;
      pdl25     : out std_logic;
      l25       : in  std_logic;
      pdl24     : out std_logic;
      l24       : in  std_logic;
      pdl23     : out std_logic;
      l23       : in  std_logic;
      pdl22     : out std_logic;
      l22       : in  std_logic;
      pdl17     : out std_logic;
      l17       : in  std_logic;
      pdl16     : out std_logic;
      l16       : in  std_logic
      );
  end component;

  component cadr_pdl1 is
    port (
      \-pdla0a\ : in  std_logic;
      \-pdla1a\ : in  std_logic;
      \-pdla2a\ : in  std_logic;
      \-pdla3a\ : in  std_logic;
      \-pdla4a\ : in  std_logic;
      pdl13     : out std_logic;
      \-pdla5a\ : in  std_logic;
      \-pdla6a\ : in  std_logic;
      \-pdla7a\ : in  std_logic;
      \-pdla8a\ : in  std_logic;
      \-pdla9a\ : in  std_logic;
      \-pwpb\   : in  std_logic;
      l13       : in  std_logic;
      pdl12     : out std_logic;
      l12       : in  std_logic;
      pdl11     : out std_logic;
      l11       : in  std_logic;
      pdl10     : out std_logic;
      \-pwpc\   : in  std_logic;
      l10       : in  std_logic;
      pdl4      : out std_logic;
      l4        : in  std_logic;
      pdl3      : out std_logic;
      l3        : in  std_logic;
      pdl2      : out std_logic;
      l2        : in  std_logic;
      pdl1      : out std_logic;
      l1        : in  std_logic;
      pdl0      : out std_logic;
      l0        : in  std_logic;
      pdl15     : out std_logic;
      l15       : in  std_logic;
      pdl14     : out std_logic;
      l14       : in  std_logic;
      pdl9      : out std_logic;
      l9        : in  std_logic;
      pdl8      : out std_logic;
      l8        : in  std_logic;
      pdl7      : out std_logic;
      l7        : in  std_logic;
      pdl6      : out std_logic;
      l6        : in  std_logic;
      pdl5      : out std_logic;
      l5        : in  std_logic
      );
  end component;

  component cadr_pdlctl is
    port (
      \-reset\      : in  std_logic;
      pdlwrited     : out std_logic;
      \-pdlwrited\  : out std_logic;
      pdlwrite      : out std_logic;
      \-destpdl(x)\ : in  std_logic;
      pwidx         : out std_logic;
      \-pwidx\      : out std_logic;
      clk4f         : in  std_logic;
      imodd         : out std_logic;
      \-imodd\      : out std_logic;
      imod          : in  std_logic;
      \-destspc\    : in  std_logic;
      \-destspcd\   : out std_logic;
      \-pdlpb\      : out std_logic;
      pdlptr0       : in  std_logic;
      pdlidx0       : in  std_logic;
      \-pdla0b\     : out std_logic;
      pdlptr1       : in  std_logic;
      pdlidx1       : in  std_logic;
      \-pdla1b\     : out std_logic;
      \-pdla2b\     : out std_logic;
      pdlidx2       : in  std_logic;
      pdlptr2       : in  std_logic;
      \-pdla3b\     : out std_logic;
      pdlidx3       : in  std_logic;
      pdlptr3       : in  std_logic;
      \-pdlpa\      : out std_logic;
      pdlptr8       : in  std_logic;
      pdlidx8       : in  std_logic;
      \-pdla8b\     : out std_logic;
      pdlptr9       : in  std_logic;
      pdlidx9       : in  std_logic;
      \-pdla9b\     : out std_logic;
      \-pdla0a\     : out std_logic;
      \-pdla1a\     : out std_logic;
      \-pdla2a\     : out std_logic;
      \-pdla3a\     : out std_logic;
      \-pdla4a\     : out std_logic;
      pdlidx4       : in  std_logic;
      pdlptr4       : in  std_logic;
      \-pdla5a\     : out std_logic;
      pdlidx5       : in  std_logic;
      pdlptr5       : in  std_logic;
      \-destpdl(p)\ : in  std_logic;
      \-pdlcnt\     : out std_logic;
      clk4b         : in  std_logic;
      ir30          : in  std_logic;
      \-clk4e\      : in  std_logic;
      \-srcpdlpop\  : in  std_logic;
      \-srcpdltop\  : in  std_logic;
      pdlenb        : out std_logic;
      tse4b         : in  std_logic;
      \-pdldrive\   : out std_logic;
      \-destpdltop\ : in  std_logic;
      \-pdla4b\     : out std_logic;
      \-pdla5b\     : out std_logic;
      \-pdla6b\     : out std_logic;
      pdlidx6       : in  std_logic;
      pdlptr6       : in  std_logic;
      \-pdla7b\     : out std_logic;
      pdlidx7       : in  std_logic;
      pdlptr7       : in  std_logic;
      wp4a          : in  std_logic;
      \-pwpa\       : out std_logic;
      \-pwpb\       : out std_logic;
      \-pwpc\       : out std_logic;
      \-pdla6a\     : out std_logic;
      \-pdla7a\     : out std_logic;
      \-pdla8a\     : out std_logic;
      \-pdla9a\     : out std_logic;
      nop           : in  std_logic
      );
  end component;

  component cadr_pdlptr is
    port (
      \-srcpdlpop\ : in  std_logic;
      clk3f        : in  std_logic;
      ob8          : in  std_logic;
      ob9          : in  std_logic;
      \-destpdlp\  : in  std_logic;
      \-pdlcry7\   : out std_logic;
      pdlptr9      : out std_logic;
      pdlptr8      : out std_logic;
      \-destpdlx\  : in  std_logic;
      pdlidx6      : out std_logic;
      ob6          : in  std_logic;
      ob7          : in  std_logic;
      pdlidx7      : out std_logic;
      pdlidx8      : out std_logic;
      pdlidx9      : out std_logic;
      ob4          : in  std_logic;
      ob5          : in  std_logic;
      \-pdlcry3\   : out std_logic;
      pdlptr7      : out std_logic;
      pdlptr6      : out std_logic;
      pdlptr5      : out std_logic;
      pdlptr4      : out std_logic;
      pdlidx0      : out std_logic;
      ob0          : in  std_logic;
      ob1          : in  std_logic;
      pdlidx1      : out std_logic;
      ob2          : in  std_logic;
      pdlidx2      : out std_logic;
      pdlidx3      : out std_logic;
      ob3          : in  std_logic;
      pdlidx4      : out std_logic;
      pdlidx5      : out std_logic;
      \-pdlcnt\    : in  std_logic;
      pdlptr3      : out std_logic;
      pdlptr2      : out std_logic;
      pdlptr1      : out std_logic;
      pdlptr0      : out std_logic;
      \-ppdrive\   : out std_logic;
      mf0          : out std_logic;
      mf1          : out std_logic;
      mf2          : out std_logic;
      mf3          : out std_logic;
      pidrive      : out std_logic;
      mf8          : out std_logic;
      mf9          : out std_logic;
      mf10         : out std_logic;
      mf11         : out std_logic;
      mf4          : out std_logic;
      mf5          : out std_logic;
      mf6          : out std_logic;
      mf7          : out std_logic;
      srcpdlidx    : in  std_logic;
      tse4b        : in  std_logic;
      srcpdlptr    : in  std_logic
      );
  end component;

  component cadr_platch is
    port (
      \-pdldrive\ : in  std_logic;
      m15         : out std_logic;
      pdl15       : in  std_logic;
      pdl14       : in  std_logic;
      m14         : out std_logic;
      m13         : out std_logic;
      pdl13       : in  std_logic;
      pdl12       : in  std_logic;
      m12         : out std_logic;
      clk4a       : in  std_logic;
      m11         : out std_logic;
      pdl11       : in  std_logic;
      pdl10       : in  std_logic;
      m10         : out std_logic;
      m9          : out std_logic;
      pdl9        : in  std_logic;
      pdl8        : in  std_logic;
      m8          : out std_logic;
      m7          : out std_logic;
      pdl7        : in  std_logic;
      pdl6        : in  std_logic;
      m6          : out std_logic;
      m5          : out std_logic;
      pdl5        : in  std_logic;
      pdl4        : in  std_logic;
      m4          : out std_logic;
      m3          : out std_logic;
      pdl3        : in  std_logic;
      pdl2        : in  std_logic;
      m2          : out std_logic;
      m1          : out std_logic;
      pdl1        : in  std_logic;
      pdl0        : in  std_logic;
      m0          : out std_logic;
      m31         : out std_logic;
      pdl31       : in  std_logic;
      pdl30       : in  std_logic;
      m30         : out std_logic;
      m29         : out std_logic;
      pdl29       : in  std_logic;
      pdl28       : in  std_logic;
      m28         : out std_logic;
      m27         : out std_logic;
      pdl27       : in  std_logic;
      pdl26       : in  std_logic;
      m26         : out std_logic;
      m25         : out std_logic;
      pdl25       : in  std_logic;
      pdl24       : in  std_logic;
      m24         : out std_logic;
      m23         : out std_logic;
      pdl23       : in  std_logic;
      pdl22       : in  std_logic;
      m22         : out std_logic;
      m21         : out std_logic;
      pdl21       : in  std_logic;
      pdl20       : in  std_logic;
      m20         : out std_logic;
      m19         : out std_logic;
      pdl19       : in  std_logic;
      pdl18       : in  std_logic;
      m18         : out std_logic;
      m17         : out std_logic;
      pdl17       : in  std_logic;
      pdl16       : in  std_logic;
      m16         : out std_logic;
      pdlparity   : in  std_logic;
      mparity     : out std_logic
      );
  end component;

  component cadr_q is
    port (
      q23      : out std_logic;
      alu24    : in  std_logic;
      alu25    : in  std_logic;
      alu26    : in  std_logic;
      alu27    : in  std_logic;
      q28      : out std_logic;
      qs0      : in  std_logic;
      qs1      : in  std_logic;
      clk2b    : in  std_logic;
      q27      : out std_logic;
      q26      : out std_logic;
      q25      : out std_logic;
      q24      : out std_logic;
      alu28    : in  std_logic;
      alu29    : in  std_logic;
      alu30    : in  std_logic;
      alu31    : in  std_logic;
      alu0     : in  std_logic;
      q31      : out std_logic;
      q30      : out std_logic;
      q29      : out std_logic;
      q15      : out std_logic;
      alu16    : in  std_logic;
      alu17    : in  std_logic;
      alu18    : in  std_logic;
      alu19    : in  std_logic;
      q20      : out std_logic;
      q19      : out std_logic;
      q18      : out std_logic;
      q17      : out std_logic;
      q16      : out std_logic;
      alu20    : in  std_logic;
      alu21    : in  std_logic;
      alu22    : in  std_logic;
      alu23    : in  std_logic;
      q22      : out std_logic;
      q21      : out std_logic;
      q7       : out std_logic;
      alu8     : in  std_logic;
      alu9     : in  std_logic;
      alu10    : in  std_logic;
      alu11    : in  std_logic;
      q12      : out std_logic;
      q11      : out std_logic;
      q10      : out std_logic;
      q9       : out std_logic;
      q8       : out std_logic;
      alu12    : in  std_logic;
      alu13    : in  std_logic;
      alu14    : in  std_logic;
      alu15    : in  std_logic;
      q14      : out std_logic;
      q13      : out std_logic;
      \-alu31\ : in  std_logic;
      alu1     : in  std_logic;
      alu2     : in  std_logic;
      alu3     : in  std_logic;
      q3       : out std_logic;
      q2       : out std_logic;
      q1       : out std_logic;
      q0       : out std_logic;
      alu4     : in  std_logic;
      alu5     : in  std_logic;
      alu6     : in  std_logic;
      alu7     : in  std_logic;
      q6       : out std_logic;
      q5       : out std_logic;
      q4       : out std_logic
      );
  end component;

  component cadr_qctl is
    port (
      \-qdrive\ : out std_logic;
      tse2      : in  std_logic;
      srcq      : out std_logic;
      q7        : in  std_logic;
      mf0       : out std_logic;
      q6        : in  std_logic;
      mf1       : out std_logic;
      q5        : in  std_logic;
      mf2       : out std_logic;
      q4        : in  std_logic;
      mf3       : out std_logic;
      q3        : in  std_logic;
      mf4       : out std_logic;
      q2        : in  std_logic;
      mf5       : out std_logic;
      q1        : in  std_logic;
      mf6       : out std_logic;
      q0        : in  std_logic;
      mf7       : out std_logic;
      qdrive    : out std_logic;
      q31       : in  std_logic;
      mf24      : out std_logic;
      q30       : in  std_logic;
      mf25      : out std_logic;
      q29       : in  std_logic;
      mf26      : out std_logic;
      q28       : in  std_logic;
      mf27      : out std_logic;
      q27       : in  std_logic;
      mf28      : out std_logic;
      q26       : in  std_logic;
      mf29      : out std_logic;
      q25       : in  std_logic;
      mf30      : out std_logic;
      q24       : in  std_logic;
      mf31      : out std_logic;
      q23       : in  std_logic;
      mf16      : out std_logic;
      q22       : in  std_logic;
      mf17      : out std_logic;
      q21       : in  std_logic;
      mf18      : out std_logic;
      q20       : in  std_logic;
      mf19      : out std_logic;
      q19       : in  std_logic;
      mf20      : out std_logic;
      q18       : in  std_logic;
      mf21      : out std_logic;
      q17       : in  std_logic;
      mf22      : out std_logic;
      q16       : in  std_logic;
      mf23      : out std_logic;
      q15       : in  std_logic;
      mf8       : out std_logic;
      q14       : in  std_logic;
      mf9       : out std_logic;
      q13       : in  std_logic;
      mf10      : out std_logic;
      q12       : in  std_logic;
      mf11      : out std_logic;
      q11       : in  std_logic;
      mf12      : out std_logic;
      q10       : in  std_logic;
      mf13      : out std_logic;
      q9        : in  std_logic;
      mf14      : out std_logic;
      q8        : in  std_logic;
      mf15      : out std_logic;
      \-srcq\   : in  std_logic;
      \-alu31\  : out std_logic;
      alu31     : in  std_logic;
      \-iralu\  : in  std_logic;
      \-ir1\    : in  std_logic;
      qs1       : out std_logic;
      \-ir0\    : in  std_logic;
      qs0       : out std_logic
      );
  end component;

  component cadr_shift0 is
    port (
      m5    : out std_logic;
      m6    : in  std_logic;
      m7    : in  std_logic;
      m8    : in  std_logic;
      m9    : in  std_logic;
      m10   : in  std_logic;
      m11   : in  std_logic;
      s1    : in  std_logic;
      s0    : in  std_logic;
      sa11  : out std_logic;
      sa10  : out std_logic;
      sa9   : out std_logic;
      sa8   : out std_logic;
      m29   : in  std_logic;
      m30   : in  std_logic;
      m31   : in  std_logic;
      m0    : in  std_logic;
      m1    : in  std_logic;
      m2    : in  std_logic;
      m3    : in  std_logic;
      sa3   : out std_logic;
      sa2   : out std_logic;
      sa1   : out std_logic;
      sa0   : out std_logic;
      m12   : in  std_logic;
      m13   : in  std_logic;
      m14   : in  std_logic;
      m15   : in  std_logic;
      sa15  : out std_logic;
      sa14  : out std_logic;
      sa12  : out std_logic;
      m4    : in  std_logic;
      sa7   : out std_logic;
      sa6   : out std_logic;
      sa5   : out std_logic;
      sa4   : out std_logic;
      sa18  : in  std_logic;
      sa22  : in  std_logic;
      sa26  : in  std_logic;
      sa30  : in  std_logic;
      s3a   : in  std_logic;
      s2a   : in  std_logic;
      r14   : out std_logic;
      r10   : out std_logic;
      \-s4\ : in  std_logic;
      r6    : out std_logic;
      r2    : out std_logic;
      s4    : in  std_logic;
      sa19  : in  std_logic;
      sa23  : in  std_logic;
      sa27  : in  std_logic;
      sa31  : in  std_logic;
      r15   : out std_logic;
      r11   : out std_logic;
      r7    : out std_logic;
      r3    : out std_logic;
      sa16  : in  std_logic;
      sa20  : in  std_logic;
      sa24  : in  std_logic;
      sa28  : in  std_logic;
      r12   : out std_logic;
      r8    : out std_logic;
      r4    : out std_logic;
      r0    : out std_logic;
      sa17  : in  std_logic;
      sa21  : in  std_logic;
      sa25  : in  std_logic;
      sa29  : in  std_logic;
      r13   : out std_logic;
      r9    : out std_logic;
      r5    : out std_logic;
      r1    : out std_logic;
      sa13  : out std_logic
      );
  end component;

  component cadr_shift1 is
    port (
      m21   : in  std_logic;
      m22   : in  std_logic;
      m23   : in  std_logic;
      m24   : in  std_logic;
      m25   : in  std_logic;
      m26   : in  std_logic;
      m27   : in  std_logic;
      s1    : in  std_logic;
      s0    : in  std_logic;
      sa27  : out std_logic;
      sa26  : out std_logic;
      sa25  : out std_logic;
      sa24  : out std_logic;
      m13   : in  std_logic;
      m14   : in  std_logic;
      m15   : in  std_logic;
      m16   : in  std_logic;
      m17   : in  std_logic;
      m18   : in  std_logic;
      m19   : in  std_logic;
      sa19  : out std_logic;
      sa18  : out std_logic;
      sa17  : out std_logic;
      sa16  : out std_logic;
      m28   : in  std_logic;
      m29   : in  std_logic;
      m30   : in  std_logic;
      m31   : in  std_logic;
      sa31  : out std_logic;
      sa30  : out std_logic;
      sa28  : out std_logic;
      m20   : in  std_logic;
      sa23  : out std_logic;
      sa22  : out std_logic;
      sa21  : out std_logic;
      sa20  : out std_logic;
      sa2   : in  std_logic;
      sa6   : in  std_logic;
      sa10  : in  std_logic;
      sa14  : in  std_logic;
      s3b   : in  std_logic;
      s2b   : in  std_logic;
      r30   : out std_logic;
      r26   : out std_logic;
      \-s4\ : in  std_logic;
      r22   : out std_logic;
      r18   : out std_logic;
      s4    : in  std_logic;
      sa3   : in  std_logic;
      sa7   : in  std_logic;
      sa11  : in  std_logic;
      sa15  : in  std_logic;
      r31   : out std_logic;
      r27   : out std_logic;
      r23   : out std_logic;
      r19   : out std_logic;
      sa0   : in  std_logic;
      sa4   : in  std_logic;
      sa8   : in  std_logic;
      sa12  : in  std_logic;
      r28   : out std_logic;
      r24   : out std_logic;
      r20   : out std_logic;
      r16   : out std_logic;
      sa1   : in  std_logic;
      sa5   : in  std_logic;
      sa9   : in  std_logic;
      sa13  : in  std_logic;
      r29   : out std_logic;
      r25   : out std_logic;
      r21   : out std_logic;
      r17   : out std_logic;
      sa29  : out std_logic
      );
  end component;

  component cadr_smctl is
    port (
      \-sr\     : out std_logic;
      \-s4\     : out std_logic;
      \-mr\     : out std_logic;
      \-irbyte\ : in  std_logic;
      ir13      : in  std_logic;
      ir12      : in  std_logic;
      \-ir0\    : in  std_logic;
      s0        : out std_logic;
      \-ir1\    : in  std_logic;
      s1        : out std_logic;
      mskl4     : out std_logic;
      ir9       : in  std_logic;
      mskr4     : out std_logic;
      mskl3cry  : out std_logic;
      s3a       : out std_logic;
      \-sh3\    : in  std_logic;
      s3b       : out std_logic;
      \-ir2\    : in  std_logic;
      s2a       : out std_logic;
      s2b       : out std_logic;
      s4        : out std_logic;
      mskr0     : out std_logic;
      mskr1     : out std_logic;
      mskr2     : out std_logic;
      mskl1     : out std_logic;
      ir6       : in  std_logic;
      mskl0     : out std_logic;
      ir5       : in  std_logic;
      mskl3     : out std_logic;
      mskr3     : out std_logic;
      ir8       : in  std_logic;
      mskl2     : out std_logic;
      ir7       : in  std_logic;
      \-sh4\    : in  std_logic
      );
  end component;

  component cadr_source is
    port (
      \-iralu\      : out std_logic;
      \-irbyte\     : out std_logic;
      dest          : out std_logic;
      \-destmem\    : out std_logic;
      ir23          : in  std_logic;
      destm         : out std_logic;
      \-specalu\    : out std_logic;
      ir8           : in  std_logic;
      iralu         : out std_logic;
      ir22          : in  std_logic;
      \-ir22\       : out std_logic;
      ir25          : in  std_logic;
      \-ir25\       : out std_logic;
      irdisp        : out std_logic;
      \-irdisp\     : out std_logic;
      irjump        : out std_logic;
      \-irjump\     : out std_logic;
      ir3           : in  std_logic;
      ir4           : in  std_logic;
      \-mul\        : out std_logic;
      \-div\        : out std_logic;
      nop           : in  std_logic;
      ir43          : in  std_logic;
      ir44          : in  std_logic;
      \-funct3\     : out std_logic;
      \-funct2\     : out std_logic;
      \-funct1\     : out std_logic;
      \-funct0\     : out std_logic;
      ir11          : in  std_logic;
      ir10          : in  std_logic;
      ir19          : in  std_logic;
      ir20          : in  std_logic;
      ir21          : in  std_logic;
      \-destintctl\ : out std_logic;
      \-destlc\     : out std_logic;
      \-destimod1\  : out std_logic;
      \-destimod0\  : out std_logic;
      \-destspc\    : out std_logic;
      \-destpdlp\   : out std_logic;
      \-destpdlx\   : out std_logic;
      \-destpdl(x)\ : out std_logic;
      \-destpdl(p)\ : out std_logic;
      \-destpdltop\ : out std_logic;
      ir26          : in  std_logic;
      ir27          : in  std_logic;
      ir28          : in  std_logic;
      \-ir31\       : in  std_logic;
      ir29          : in  std_logic;
      \-srcq\       : out std_logic;
      \-srcopc\     : out std_logic;
      \-srcpdltop\  : out std_logic;
      \-srcpdlpop\  : out std_logic;
      \-srcpdlidx\  : out std_logic;
      \-srcpdlptr\  : out std_logic;
      \-srcspc\     : out std_logic;
      \-srcdc\      : out std_logic;
      \-srcspcpop\  : out std_logic;
      \-srclc\      : out std_logic;
      \-srcmd\      : out std_logic;
      \-srcmap\     : out std_logic;
      \-srcvma\     : out std_logic;
      \destimod0 l\ : in  std_logic;
      \iwrited l\   : in  std_logic;
      \-destmdr\    : out std_logic;
      \-destvma\    : out std_logic;
      \-idebug\     : in  std_logic;
      imod          : out std_logic
      );
  end component;

  component cadr_spc is
    port (
      \-swpa\   : in  std_logic;
      spcw14    : in  std_logic;
      spcptr4   : out std_logic;
      spco14    : out std_logic;
      spco15    : out std_logic;
      spcptr3   : out std_logic;
      spcptr2   : out std_logic;
      spcptr1   : out std_logic;
      spcptr0   : out std_logic;
      spcw15    : in  std_logic;
      spcw12    : in  std_logic;
      spco12    : out std_logic;
      spco13    : out std_logic;
      spcw13    : in  std_logic;
      spcw10    : in  std_logic;
      spco10    : out std_logic;
      spco11    : out std_logic;
      spcw11    : in  std_logic;
      spcopar   : out std_logic;
      spco18    : out std_logic;
      spco17    : out std_logic;
      spco16    : out std_logic;
      \-swpb\   : in  std_logic;
      spcw4     : in  std_logic;
      spco4     : out std_logic;
      spco5     : out std_logic;
      spcw5     : in  std_logic;
      spcw2     : in  std_logic;
      spco2     : out std_logic;
      spco3     : out std_logic;
      spcw3     : in  std_logic;
      spcw0     : in  std_logic;
      spco0     : out std_logic;
      spco1     : out std_logic;
      spcw1     : in  std_logic;
      spco9     : out std_logic;
      spco8     : out std_logic;
      spco7     : out std_logic;
      spco6     : out std_logic;
      spush     : in  std_logic;
      clk4f     : in  std_logic;
      \-spcnt\  : in  std_logic;
      \-spccry\ : out std_logic;
      spcw18    : in  std_logic;
      spcwpar   : in  std_logic;
      spcw16    : in  std_logic;
      spcw17    : in  std_logic;
      spcw8     : in  std_logic;
      spcw9     : in  std_logic;
      spcw6     : in  std_logic;
      spcw7     : in  std_logic
      );
  end component;

  component cadr_spclch is
    port (
      \-spcdrive\ : in  std_logic;
      m23         : out std_logic;
      m22         : out std_logic;
      m21         : out std_logic;
      m20         : out std_logic;
      clk4c       : in  std_logic;
      m19         : out std_logic;
      spco18      : in  std_logic;
      m18         : out std_logic;
      m17         : out std_logic;
      spco17      : in  std_logic;
      spco16      : in  std_logic;
      m16         : out std_logic;
      m15         : out std_logic;
      spco15      : in  std_logic;
      spco14      : in  std_logic;
      m14         : out std_logic;
      m13         : out std_logic;
      spco13      : in  std_logic;
      spco12      : in  std_logic;
      m12         : out std_logic;
      m11         : out std_logic;
      spco11      : in  std_logic;
      spco10      : in  std_logic;
      m10         : out std_logic;
      m9          : out std_logic;
      spco9       : in  std_logic;
      spco8       : in  std_logic;
      m8          : out std_logic;
      m7          : out std_logic;
      spco7       : in  std_logic;
      spco6       : in  std_logic;
      m6          : out std_logic;
      m5          : out std_logic;
      spco5       : in  std_logic;
      spco4       : in  std_logic;
      m4          : out std_logic;
      m3          : out std_logic;
      spco3       : in  std_logic;
      spco2       : in  std_logic;
      m2          : out std_logic;
      m1          : out std_logic;
      spco1       : in  std_logic;
      spco0       : in  std_logic;
      m0          : out std_logic;
      m24         : out std_logic;
      m25         : out std_logic;
      m26         : out std_logic;
      spcptr4     : in  std_logic;
      m27         : out std_logic;
      spcptr3     : in  std_logic;
      m28         : out std_logic;
      spcptr2     : in  std_logic;
      m29         : out std_logic;
      spcptr1     : in  std_logic;
      m30         : out std_logic;
      spcptr0     : in  std_logic;
      m31         : out std_logic;
      spcdrive    : in  std_logic;
      spc16       : out std_logic;
      spc17       : out std_logic;
      spc18       : out std_logic;
      spcpar      : out std_logic;
      spcwpar     : in  std_logic;
      spcw18      : in  std_logic;
      spcw17      : in  std_logic;
      spcw16      : in  std_logic;
      spcwpass    : in  std_logic;
      \-spcwpass\ : in  std_logic;
      spcw15      : in  std_logic;
      spc8        : out std_logic;
      spcw14      : in  std_logic;
      spc9        : out std_logic;
      spcw13      : in  std_logic;
      spc10       : out std_logic;
      spcw12      : in  std_logic;
      spc11       : out std_logic;
      spcw11      : in  std_logic;
      spc12       : out std_logic;
      spcw10      : in  std_logic;
      spc13       : out std_logic;
      spcw9       : in  std_logic;
      spc14       : out std_logic;
      spcw8       : in  std_logic;
      spc15       : out std_logic;
      spcw7       : in  std_logic;
      spcw6       : in  std_logic;
      spc1        : out std_logic;
      spcw5       : in  std_logic;
      spc2        : out std_logic;
      spcw4       : in  std_logic;
      spc3        : out std_logic;
      spcw3       : in  std_logic;
      spc4        : out std_logic;
      spcw2       : in  std_logic;
      spc5        : out std_logic;
      spcw1       : in  std_logic;
      spc6        : out std_logic;
      spcw0       : in  std_logic;
      spc7        : out std_logic;
      \-spcpass\  : in  std_logic;
      clk4d       : in  std_logic;
      spcopar     : in  std_logic;
      spc0        : out std_logic
      );
  end component;

  component cadr_spcpar is
    port (
      spcwparh    : out std_logic;
      \-spcwparl\ : out std_logic;
      spcwpar     : out std_logic;
      spcw17      : in  std_logic;
      spcw18      : in  std_logic;
      spcw12      : in  std_logic;
      spcw13      : in  std_logic;
      spcw14      : in  std_logic;
      spcw15      : in  std_logic;
      spcw16      : in  std_logic;
      spcw5       : in  std_logic;
      spcw6       : in  std_logic;
      spcw7       : in  std_logic;
      spcw8       : in  std_logic;
      spcw9       : in  std_logic;
      spcw10      : in  std_logic;
      spcw11      : in  std_logic;
      spcw0       : in  std_logic;
      spcw1       : in  std_logic;
      spcw2       : in  std_logic;
      spcw3       : in  std_logic;
      spcw4       : in  std_logic;
      spc16       : in  std_logic;
      spc17       : in  std_logic;
      spc18       : in  std_logic;
      spcpar      : in  std_logic;
      spcparh     : out std_logic;
      spc11       : in  std_logic;
      spc12       : in  std_logic;
      spc13       : in  std_logic;
      spc14       : in  std_logic;
      spc15       : in  std_logic;
      spc5        : in  std_logic;
      spc6        : in  std_logic;
      spc7        : in  std_logic;
      spc8        : in  std_logic;
      spc9        : in  std_logic;
      spc10       : in  std_logic;
      spcparok    : out std_logic;
      spc0        : in  std_logic;
      spc1        : in  std_logic;
      spc2        : in  std_logic;
      spc3        : in  std_logic;
      spc4        : in  std_logic
      );
  end component;

  component cadr_spcw is
    port (
      destspcd : in  std_logic;
      reta12   : out std_logic;
      l12      : in  std_logic;
      spcw12   : out std_logic;
      reta13   : out std_logic;
      l13      : in  std_logic;
      spcw13   : out std_logic;
      spcw14   : out std_logic;
      l14      : in  std_logic;
      spcw15   : out std_logic;
      l15      : in  std_logic;
      reta8    : out std_logic;
      l8       : in  std_logic;
      spcw8    : out std_logic;
      reta9    : out std_logic;
      l9       : in  std_logic;
      spcw9    : out std_logic;
      spcw10   : out std_logic;
      l10      : in  std_logic;
      reta10   : out std_logic;
      spcw11   : out std_logic;
      l11      : in  std_logic;
      reta11   : out std_logic;
      reta4    : out std_logic;
      l4       : in  std_logic;
      spcw4    : out std_logic;
      reta5    : out std_logic;
      l5       : in  std_logic;
      spcw5    : out std_logic;
      spcw6    : out std_logic;
      l6       : in  std_logic;
      reta6    : out std_logic;
      spcw7    : out std_logic;
      l7       : in  std_logic;
      reta7    : out std_logic;
      reta0    : out std_logic;
      l0       : in  std_logic;
      spcw0    : out std_logic;
      reta1    : out std_logic;
      l1       : in  std_logic;
      spcw1    : out std_logic;
      spcw2    : out std_logic;
      l2       : in  std_logic;
      reta2    : out std_logic;
      spcw3    : out std_logic;
      l3       : in  std_logic;
      reta3    : out std_logic;
      n        : in  std_logic;
      ipc12    : in  std_logic;
      wpc12    : in  std_logic;
      wpc13    : in  std_logic;
      ipc13    : in  std_logic;
      clk4d    : in  std_logic;
      ipc8     : in  std_logic;
      wpc8     : in  std_logic;
      wpc9     : in  std_logic;
      ipc9     : in  std_logic;
      ipc10    : in  std_logic;
      wpc10    : in  std_logic;
      wpc11    : in  std_logic;
      ipc11    : in  std_logic;
      ipc4     : in  std_logic;
      wpc4     : in  std_logic;
      wpc5     : in  std_logic;
      ipc5     : in  std_logic;
      ipc6     : in  std_logic;
      wpc6     : in  std_logic;
      wpc7     : in  std_logic;
      ipc7     : in  std_logic;
      ipc0     : in  std_logic;
      wpc0     : in  std_logic;
      wpc1     : in  std_logic;
      ipc1     : in  std_logic;
      ipc2     : in  std_logic;
      wpc2     : in  std_logic;
      wpc3     : in  std_logic;
      ipc3     : in  std_logic;
      l16      : in  std_logic;
      spcw16   : out std_logic;
      l17      : in  std_logic;
      spcw17   : out std_logic;
      spcw18   : out std_logic;
      l18      : in  std_logic
      );
  end component;

  component cadr_spy1 is
    port (
      \-spy.obl\ : out std_logic;
      ob7        : in  std_logic;
      spy0       : out std_logic;
      ob6        : in  std_logic;
      spy1       : out std_logic;
      ob5        : in  std_logic;
      spy2       : out std_logic;
      ob4        : in  std_logic;
      spy3       : out std_logic;
      ob3        : in  std_logic;
      spy4       : out std_logic;
      ob2        : in  std_logic;
      spy5       : out std_logic;
      ob1        : in  std_logic;
      spy6       : out std_logic;
      ob0        : in  std_logic;
      spy7       : out std_logic;
      ob15       : in  std_logic;
      spy8       : out std_logic;
      ob14       : in  std_logic;
      spy9       : out std_logic;
      ob13       : in  std_logic;
      spy10      : out std_logic;
      ob12       : in  std_logic;
      spy11      : out std_logic;
      ob11       : in  std_logic;
      spy12      : out std_logic;
      ob10       : in  std_logic;
      spy13      : out std_logic;
      ob9        : in  std_logic;
      spy14      : out std_logic;
      ob8        : in  std_logic;
      spy15      : out std_logic;
      \-spy.obh\ : in  std_logic;
      ob23       : in  std_logic;
      ob22       : in  std_logic;
      ob21       : in  std_logic;
      ob20       : in  std_logic;
      ob19       : in  std_logic;
      ob18       : in  std_logic;
      ob17       : in  std_logic;
      ob16       : in  std_logic;
      ob31       : in  std_logic;
      ob30       : in  std_logic;
      ob29       : in  std_logic;
      ob28       : in  std_logic;
      ob27       : in  std_logic;
      ob26       : in  std_logic;
      ob25       : in  std_logic;
      ob24       : in  std_logic;
      \-spy.irl\ : in  std_logic;
      ir7        : in  std_logic;
      ir6        : in  std_logic;
      ir5        : in  std_logic;
      ir4        : in  std_logic;
      ir3        : in  std_logic;
      ir2        : in  std_logic;
      ir1        : in  std_logic;
      ir0        : in  std_logic;
      ir15       : in  std_logic;
      ir14       : in  std_logic;
      ir13       : in  std_logic;
      ir12       : in  std_logic;
      ir11       : in  std_logic;
      ir10       : in  std_logic;
      ir9        : in  std_logic;
      ir8        : in  std_logic;
      \-spy.irh\ : in  std_logic;
      ir47       : in  std_logic;
      ir46       : in  std_logic;
      ir45       : in  std_logic;
      ir44       : in  std_logic;
      ir43       : in  std_logic;
      ir42       : in  std_logic;
      ir41       : in  std_logic;
      ir40       : in  std_logic;
      ir39       : in  std_logic;
      ir38       : in  std_logic;
      ir37       : in  std_logic;
      ir36       : in  std_logic;
      ir35       : in  std_logic;
      ir34       : in  std_logic;
      ir33       : in  std_logic;
      ir32       : in  std_logic;
      \-spy.irm\ : in  std_logic;
      ir31       : in  std_logic;
      ir30       : in  std_logic;
      ir29       : in  std_logic;
      ir28       : in  std_logic;
      ir27       : in  std_logic;
      ir26       : in  std_logic;
      ir25       : in  std_logic;
      ir24       : in  std_logic;
      ir23       : in  std_logic;
      ir22       : in  std_logic;
      ir21       : in  std_logic;
      ir20       : in  std_logic;
      ir19       : in  std_logic;
      ir18       : in  std_logic;
      ir17       : in  std_logic;
      ir16       : in  std_logic
      );
  end component;

  component cadr_spy2 is
    port (
      \-spy.al\    : out std_logic;
      aa15         : in  std_logic;
      spy8         : out std_logic;
      aa14         : in  std_logic;
      spy9         : out std_logic;
      aa13         : in  std_logic;
      spy10        : out std_logic;
      aa12         : in  std_logic;
      spy11        : out std_logic;
      aa11         : in  std_logic;
      spy12        : out std_logic;
      aa10         : in  std_logic;
      spy13        : out std_logic;
      aa9          : in  std_logic;
      spy14        : out std_logic;
      aa8          : in  std_logic;
      spy15        : out std_logic;
      aa7          : in  std_logic;
      spy0         : out std_logic;
      aa6          : in  std_logic;
      spy1         : out std_logic;
      aa5          : in  std_logic;
      spy2         : out std_logic;
      aa4          : in  std_logic;
      spy3         : out std_logic;
      aa3          : in  std_logic;
      spy4         : out std_logic;
      aa2          : in  std_logic;
      spy5         : out std_logic;
      aa1          : in  std_logic;
      spy6         : out std_logic;
      aa0          : in  std_logic;
      spy7         : out std_logic;
      \-spy.ah\    : in  std_logic;
      a31a         : in  std_logic;
      a30          : in  std_logic;
      a29          : in  std_logic;
      a28          : in  std_logic;
      a27          : in  std_logic;
      a26          : in  std_logic;
      a25          : in  std_logic;
      a24          : in  std_logic;
      a23          : in  std_logic;
      a22          : in  std_logic;
      a21          : in  std_logic;
      a20          : in  std_logic;
      a19          : in  std_logic;
      a18          : in  std_logic;
      a17          : in  std_logic;
      a16          : in  std_logic;
      \-spy.flag2\ : in  std_logic;
      ir48         : in  std_logic;
      nop          : in  std_logic;
      \-vmaok\     : in  std_logic;
      jcond        : in  std_logic;
      pcs1         : in  std_logic;
      pcs0         : in  std_logic;
      wmapd        : in  std_logic;
      destspcd     : in  std_logic;
      iwrited      : in  std_logic;
      imodd        : in  std_logic;
      pdlwrited    : in  std_logic;
      spushd       : in  std_logic;
      \-spy.ml\    : in  std_logic;
      m15          : in  std_logic;
      m14          : in  std_logic;
      m13          : in  std_logic;
      m12          : in  std_logic;
      m11          : in  std_logic;
      m10          : in  std_logic;
      m9           : in  std_logic;
      m8           : in  std_logic;
      m7           : in  std_logic;
      m6           : in  std_logic;
      m5           : in  std_logic;
      m4           : in  std_logic;
      m3           : in  std_logic;
      m2           : in  std_logic;
      m1           : in  std_logic;
      m0           : in  std_logic;
      \-spy.mh\    : in  std_logic;
      m23          : in  std_logic;
      m22          : in  std_logic;
      m21          : in  std_logic;
      m20          : in  std_logic;
      m19          : in  std_logic;
      m18          : in  std_logic;
      m17          : in  std_logic;
      m16          : in  std_logic;
      m31          : in  std_logic;
      m30          : in  std_logic;
      m29          : in  std_logic;
      m28          : in  std_logic;
      m27          : in  std_logic;
      m26          : in  std_logic;
      m25          : in  std_logic;
      m24          : in  std_logic
      );
  end component;

  component cadr_trap is
    port (
      mdparerr    : out std_logic;
      mdpareven   : out std_logic;
      mdpar       : in  std_logic;
      \-md5\      : in  std_logic;
      \-md6\      : in  std_logic;
      \-md7\      : in  std_logic;
      \-md8\      : in  std_logic;
      \-md9\      : in  std_logic;
      \-md10\     : in  std_logic;
      \-md11\     : in  std_logic;
      mdparl      : out std_logic;
      \-md0\      : in  std_logic;
      \-md1\      : in  std_logic;
      \-md2\      : in  std_logic;
      \-md3\      : in  std_logic;
      \-md4\      : in  std_logic;
      \-md17\     : in  std_logic;
      \-md18\     : in  std_logic;
      \-md19\     : in  std_logic;
      \-md20\     : in  std_logic;
      \-md21\     : in  std_logic;
      \-md22\     : in  std_logic;
      \-md23\     : in  std_logic;
      mdparm      : out std_logic;
      \-md12\     : in  std_logic;
      \-md13\     : in  std_logic;
      \-md14\     : in  std_logic;
      \-md15\     : in  std_logic;
      \-md16\     : in  std_logic;
      \-md29\     : in  std_logic;
      \-md30\     : in  std_logic;
      \-md31\     : in  std_logic;
      mdparodd    : out std_logic;
      \-md24\     : in  std_logic;
      \-md25\     : in  std_logic;
      \-md26\     : in  std_logic;
      \-md27\     : in  std_logic;
      \-md28\     : in  std_logic;
      mdhaspar    : in  std_logic;
      \use.md\    : in  std_logic;
      \-wait\     : in  std_logic;
      \-parerr\   : out std_logic;
      \-trap\     : out std_logic;
      \boot.trap\ : in  std_logic;
      \-trapenb\  : out std_logic;
      \-memparok\ : out std_logic;
      trapb       : out std_logic;
      trapa       : out std_logic;
      memparok    : out std_logic;
      trapenb     : in  std_logic
      );
  end component;

  component cadr_vctl1 is
    port (
      \-reset\             : in  std_logic;
      rdcyc                : out std_logic;
      wrcyc                : out std_logic;
      clk2a                : in  std_logic;
      wmap                 : in  std_logic;
      \-wmapd\             : out std_logic;
      wmapd                : out std_logic;
      memprepare           : out std_logic;
      \-memwr\             : in  std_logic;
      \-memprepare\        : in  std_logic;
      \-lvmo22\            : in  std_logic;
      \-pfw\               : out std_logic;
      \-pfr\               : in  std_logic;
      \-vmaok\             : out std_logic;
      \-mfinishd\          : out std_logic;
      memrq                : out std_logic;
      mclk1a               : in  std_logic;
      mbusy                : out std_logic;
      \rd.in.progress\     : out std_logic;
      \set.rd.in.progress\ : out std_logic;
      \-rdfinish\          : out std_logic;
      \-mfinish\           : out std_logic;
      clk2c                : in  std_logic;
      \-memop\             : out std_logic;
      \-memack\            : in  std_logic;
      \-memrd\             : in  std_logic;
      \-ifetch\            : in  std_logic;
      memstart             : out std_logic;
      \-memstart\          : out std_logic;
      \-mbusy.sync\        : out std_logic;
      \mbusy.sync\         : out std_logic;
      destmem              : in  std_logic;
      \-memgrant\          : in  std_logic;
      \use.md\             : in  std_logic;
      \-wait\              : out std_logic;
      needfetch            : in  std_logic;
      lcinc                : in  std_logic;
      \-hang\              : out std_logic;
      \-clk3g\             : in  std_logic
      );
  end component;

  component cadr_vctl2 is
    port (
      mapwr0d        : out std_logic;
      \-wmapd\       : out std_logic;
      \-vma26\       : in  std_logic;
      mapwr1d        : out std_logic;
      \-vma25\       : in  std_logic;
      wp1a           : in  std_logic;
      \-vm0wpa\      : out std_logic;
      \-vm0wpb\      : out std_logic;
      \-vm1wpa\      : out std_logic;
      wp1b           : in  std_logic;
      \-vm1wpb\      : out std_logic;
      \-lvmo23\      : in  std_logic;
      \-pfr\         : out std_logic;
      \-wmap\        : out std_logic;
      wmap           : out std_logic;
      \-memrq\       : out std_logic;
      memrq          : in  std_logic;
      \-memprepare\  : out std_logic;
      memprepare     : in  std_logic;
      destmem        : out std_logic;
      \-destmem\     : in  std_logic;
      mdsela         : out std_logic;
      \-destmdr\     : in  std_logic;
      clk2c          : in  std_logic;
      mdselb         : out std_logic;
      \-destvma\     : in  std_logic;
      \-ifetch\      : in  std_logic;
      \-vmaenb\      : out std_logic;
      vmasela        : out std_logic;
      vmaselb        : out std_logic;
      wrcyc          : in  std_logic;
      \lm drive enb\ : in  std_logic;
      \-memdrive.a\  : out std_logic;
      \-memdrive.b\  : out std_logic;
      \-memwr\       : out std_logic;
      \-memrd\       : out std_logic;
      ir20           : in  std_logic;
      ir19           : in  std_logic;
      \use.md\       : out std_logic;
      \-srcmd\       : in  std_logic;
      nopa           : out std_logic;
      \-nopa\        : in  std_logic
      );
  end component;

  component cadr_vma is
    port (
      \-vmadrive\ : out std_logic;
      \-vma31\    : out std_logic;
      mf24        : out std_logic;
      \-vma30\    : out std_logic;
      mf25        : out std_logic;
      \-vma29\    : out std_logic;
      mf26        : out std_logic;
      \-vma28\    : out std_logic;
      mf27        : out std_logic;
      \-vma27\    : out std_logic;
      mf28        : out std_logic;
      \-vma26\    : out std_logic;
      mf29        : out std_logic;
      \-vma25\    : out std_logic;
      mf30        : out std_logic;
      \-vma24\    : out std_logic;
      mf31        : out std_logic;
      \-vma7\     : out std_logic;
      mf0         : out std_logic;
      \-vma6\     : out std_logic;
      mf1         : out std_logic;
      \-vma5\     : out std_logic;
      mf2         : out std_logic;
      \-vma4\     : out std_logic;
      mf3         : out std_logic;
      \-vma3\     : out std_logic;
      mf4         : out std_logic;
      \-vma2\     : out std_logic;
      mf5         : out std_logic;
      \-vma1\     : out std_logic;
      mf6         : out std_logic;
      \-vma0\     : out std_logic;
      mf7         : out std_logic;
      \-vma23\    : out std_logic;
      mf16        : out std_logic;
      \-vma22\    : out std_logic;
      mf17        : out std_logic;
      \-vma21\    : out std_logic;
      mf18        : out std_logic;
      \-vma20\    : out std_logic;
      mf19        : out std_logic;
      \-vma19\    : out std_logic;
      mf20        : out std_logic;
      \-vma18\    : out std_logic;
      mf21        : out std_logic;
      \-vma17\    : out std_logic;
      mf22        : out std_logic;
      \-vma16\    : out std_logic;
      mf23        : out std_logic;
      \-vma15\    : out std_logic;
      mf8         : out std_logic;
      \-vma14\    : out std_logic;
      mf9         : out std_logic;
      \-vma13\    : out std_logic;
      mf10        : out std_logic;
      \-vma12\    : out std_logic;
      mf11        : out std_logic;
      \-vma11\    : out std_logic;
      mf12        : out std_logic;
      \-vma10\    : out std_logic;
      mf13        : out std_logic;
      \-vma9\     : out std_logic;
      mf14        : out std_logic;
      \-vma8\     : out std_logic;
      mf15        : out std_logic;
      tse2        : in  std_logic;
      \-vmaenb\   : in  std_logic;
      \-vmas24\   : in  std_logic;
      \-vmas25\   : in  std_logic;
      \-vmas26\   : in  std_logic;
      clk1a       : in  std_logic;
      \-vmas27\   : in  std_logic;
      \-vmas28\   : in  std_logic;
      \-vmas29\   : in  std_logic;
      \-vmas30\   : in  std_logic;
      \-vmas31\   : in  std_logic;
      \-vmas0\    : in  std_logic;
      \-vmas1\    : in  std_logic;
      \-vmas2\    : in  std_logic;
      clk2a       : in  std_logic;
      \-vmas3\    : in  std_logic;
      \-vmas4\    : in  std_logic;
      \-vmas5\    : in  std_logic;
      \-vmas12\   : in  std_logic;
      \-vmas13\   : in  std_logic;
      \-vmas14\   : in  std_logic;
      \-vmas15\   : in  std_logic;
      \-vmas16\   : in  std_logic;
      \-vmas17\   : in  std_logic;
      \-vmas18\   : in  std_logic;
      \-vmas19\   : in  std_logic;
      \-vmas20\   : in  std_logic;
      \-vmas21\   : in  std_logic;
      \-vmas22\   : in  std_logic;
      \-vmas23\   : in  std_logic;
      \-vmas6\    : in  std_logic;
      \-vmas7\    : in  std_logic;
      \-vmas8\    : in  std_logic;
      clk2c       : in  std_logic;
      \-vmas9\    : in  std_logic;
      \-vmas10\   : in  std_logic;
      \-vmas11\   : in  std_logic;
      \-srcvma\   : in  std_logic;
      srcvma      : out std_logic
      );
  end component;

  component cadr_vmas is
    port (
      vmasela     : in  std_logic;
      lc22        : in  std_logic;
      ob20        : in  std_logic;
      \-vmas20\   : out std_logic;
      lc23        : in  std_logic;
      ob21        : in  std_logic;
      \-vmas21\   : out std_logic;
      \-vmas22\   : out std_logic;
      ob22        : in  std_logic;
      lc24        : in  std_logic;
      \-vmas23\   : out std_logic;
      ob23        : in  std_logic;
      lc25        : in  std_logic;
      ob28        : in  std_logic;
      \-vmas28\   : out std_logic;
      ob29        : in  std_logic;
      \-vmas29\   : out std_logic;
      \-vmas30\   : out std_logic;
      ob30        : in  std_logic;
      \-vmas31\   : out std_logic;
      ob31        : in  std_logic;
      vmaselb     : in  std_logic;
      lc14        : in  std_logic;
      ob12        : in  std_logic;
      \-vmas12\   : out std_logic;
      lc15        : in  std_logic;
      ob13        : in  std_logic;
      \-vmas13\   : out std_logic;
      \-vmas14\   : out std_logic;
      ob14        : in  std_logic;
      lc16        : in  std_logic;
      \-vmas15\   : out std_logic;
      ob15        : in  std_logic;
      lc17        : in  std_logic;
      lc18        : in  std_logic;
      ob16        : in  std_logic;
      \-vmas16\   : out std_logic;
      lc19        : in  std_logic;
      ob17        : in  std_logic;
      \-vmas17\   : out std_logic;
      \-vmas18\   : out std_logic;
      ob18        : in  std_logic;
      lc20        : in  std_logic;
      \-vmas19\   : out std_logic;
      ob19        : in  std_logic;
      lc21        : in  std_logic;
      \-memstart\ : in  std_logic;
      \-vma12\    : in  std_logic;
      \-md12\     : in  std_logic;
      mapi12      : out std_logic;
      \-vma13\    : in  std_logic;
      \-md13\     : in  std_logic;
      mapi13      : out std_logic;
      mapi14      : out std_logic;
      \-md14\     : in  std_logic;
      \-vma14\    : in  std_logic;
      mapi15      : out std_logic;
      \-md15\     : in  std_logic;
      \-vma15\    : in  std_logic;
      \-vma16\    : in  std_logic;
      \-md16\     : in  std_logic;
      mapi16      : out std_logic;
      \-vma17\    : in  std_logic;
      \-md17\     : in  std_logic;
      mapi17      : out std_logic;
      mapi18      : out std_logic;
      \-md18\     : in  std_logic;
      \-vma18\    : in  std_logic;
      mapi19      : out std_logic;
      \-md19\     : in  std_logic;
      \-vma19\    : in  std_logic;
      \-vma20\    : in  std_logic;
      \-md20\     : in  std_logic;
      mapi20      : out std_logic;
      \-vma21\    : in  std_logic;
      \-md21\     : in  std_logic;
      mapi21      : out std_logic;
      mapi22      : out std_logic;
      \-md22\     : in  std_logic;
      \-vma22\    : in  std_logic;
      mapi23      : out std_logic;
      \-md23\     : in  std_logic;
      \-vma23\    : in  std_logic;
      lc2         : in  std_logic;
      ob0         : in  std_logic;
      \-vmas0\    : out std_logic;
      lc3         : in  std_logic;
      ob1         : in  std_logic;
      \-vmas1\    : out std_logic;
      \-vmas2\    : out std_logic;
      ob2         : in  std_logic;
      lc4         : in  std_logic;
      \-vmas3\    : out std_logic;
      ob3         : in  std_logic;
      lc5         : in  std_logic;
      \-vma8\     : in  std_logic;
      \-md8\      : in  std_logic;
      mapi8       : out std_logic;
      \-vma9\     : in  std_logic;
      \-md9\      : in  std_logic;
      mapi9       : out std_logic;
      mapi10      : out std_logic;
      \-md10\     : in  std_logic;
      \-vma10\    : in  std_logic;
      mapi11      : out std_logic;
      \-md11\     : in  std_logic;
      \-vma11\    : in  std_logic;
      lc10        : in  std_logic;
      ob8         : in  std_logic;
      \-vmas8\    : out std_logic;
      lc11        : in  std_logic;
      ob9         : in  std_logic;
      \-vmas9\    : out std_logic;
      \-vmas10\   : out std_logic;
      ob10        : in  std_logic;
      lc12        : in  std_logic;
      \-vmas11\   : out std_logic;
      ob11        : in  std_logic;
      lc13        : in  std_logic;
      lc6         : in  std_logic;
      ob4         : in  std_logic;
      \-vmas4\    : out std_logic;
      lc7         : in  std_logic;
      ob5         : in  std_logic;
      \-vmas5\    : out std_logic;
      \-vmas6\    : out std_logic;
      ob6         : in  std_logic;
      lc8         : in  std_logic;
      \-vmas7\    : out std_logic;
      ob7         : in  std_logic;
      lc9         : in  std_logic;
      ob24        : in  std_logic;
      \-vmas24\   : out std_logic;
      ob25        : in  std_logic;
      \-vmas25\   : out std_logic;
      \-vmas26\   : out std_logic;
      ob26        : in  std_logic;
      \-vmas27\   : out std_logic;
      ob27        : in  std_logic
      );
  end component;

  component cadr_vmem0 is
    port (
      \-vmap0\   : out std_logic;
      \-vmap1\   : out std_logic;
      \-vmap2\   : out std_logic;
      \-vmap3\   : out std_logic;
      \-vmap4\   : out std_logic;
      vpari      : out std_logic;
      \-vma27\   : in  std_logic;
      \-vma28\   : in  std_logic;
      \-vma29\   : in  std_logic;
      vm0pari    : out std_logic;
      \-vma30\   : in  std_logic;
      \-vma31\   : in  std_logic;
      \-mapi23\  : out std_logic;
      mapi22     : in  std_logic;
      mapi21     : in  std_logic;
      mapi20     : in  std_logic;
      mapi19     : in  std_logic;
      mapi18     : in  std_logic;
      mapi17     : in  std_logic;
      mapi16     : in  std_logic;
      mapi15     : in  std_logic;
      mapi14     : in  std_logic;
      mapi13     : in  std_logic;
      \-vm0wpb\  : in  std_logic;
      mapi23     : in  std_logic;
      \-vm0wpa\  : in  std_logic;
      memstart   : in  std_logic;
      srcmap     : in  std_logic;
      \-use.map\ : out std_logic;
      v0parok    : out std_logic;
      vmoparodd  : in  std_logic;
      vmoparok   : out std_logic
      );
  end component;

  component cadr_vmem1 is
    port (
      \-vma17\   : in  std_logic;
      \-vma18\   : in  std_logic;
      \-vma19\   : in  std_logic;
      \-vma20\   : in  std_logic;
      \-vma21\   : in  std_logic;
      \-vma22\   : in  std_logic;
      \-vma23\   : in  std_logic;
      vm1mpar    : out std_logic;
      \-vma12\   : in  std_logic;
      \-vma13\   : in  std_logic;
      \-vma14\   : in  std_logic;
      \-vma15\   : in  std_logic;
      \-vma16\   : in  std_logic;
      \-vma5\    : in  std_logic;
      \-vma7\    : in  std_logic;
      \-vma8\    : in  std_logic;
      \-vma9\    : in  std_logic;
      \-vma10\   : in  std_logic;
      \-vma11\   : in  std_logic;
      \-vm1lpar\ : out std_logic;
      \-vma0\    : in  std_logic;
      \-vma1\    : in  std_logic;
      \-vma2\    : in  std_logic;
      \-vma3\    : in  std_logic;
      \-vma4\    : in  std_logic;
      vmap4a     : out std_logic;
      vmap3a     : out std_logic;
      vmap2a     : out std_logic;
      vmap1a     : out std_logic;
      vmap0a     : out std_logic;
      \-vmo10\   : out std_logic;
      \-mapi12a\ : out std_logic;
      \-mapi11a\ : out std_logic;
      \-mapi10a\ : out std_logic;
      \-mapi9a\  : out std_logic;
      \-mapi8a\  : out std_logic;
      \-vm1wpa\  : in  std_logic;
      \-vmo4\    : out std_logic;
      \-vmo2\    : out std_logic;
      mapi10     : in  std_logic;
      mapi9      : in  std_logic;
      mapi8      : in  std_logic;
      \-vmap4\   : in  std_logic;
      \-vmap3\   : in  std_logic;
      \-vmap2\   : in  std_logic;
      \-vmap1\   : in  std_logic;
      \-vmap0\   : in  std_logic;
      \-vmo0\    : out std_logic;
      vm1pari    : out std_logic;
      mapi12     : in  std_logic;
      mapi11     : in  std_logic;
      \-mapi8b\  : out std_logic;
      \-mapi9b\  : out std_logic;
      \-mapi10b\ : out std_logic;
      \-mapi11b\ : out std_logic;
      \-mapi12b\ : out std_logic;
      \-vmo11\   : out std_logic;
      \-vmo5\    : out std_logic;
      \-vmo9\    : out std_logic;
      \-vmo3\    : out std_logic;
      \-vmo8\    : out std_logic;
      \-vmo7\    : out std_logic;
      \-vmo1\    : out std_logic;
      \-vmo6\    : out std_logic;
      \-vma6\    : in  std_logic
      );
  end component;

  component cadr_vmem2 is
    port (
      vmap4b     : out std_logic;
      vmap3b     : out std_logic;
      vmap2b     : out std_logic;
      vmap1b     : out std_logic;
      vmap0b     : out std_logic;
      \-vmo20\   : out std_logic;
      \-mapi12b\ : in  std_logic;
      \-mapi11b\ : in  std_logic;
      \-mapi10b\ : in  std_logic;
      \-mapi9b\  : in  std_logic;
      \-mapi8b\  : in  std_logic;
      \-vm1wpb\  : in  std_logic;
      \-vma20\   : in  std_logic;
      \-vmo21\   : out std_logic;
      \-vma21\   : in  std_logic;
      \-vmo22\   : out std_logic;
      \-vma22\   : in  std_logic;
      \-vmo23\   : out std_logic;
      \-vma23\   : in  std_logic;
      \-vmo16\   : out std_logic;
      \-vma16\   : in  std_logic;
      \-vmo17\   : out std_logic;
      \-vma17\   : in  std_logic;
      \-vmo18\   : out std_logic;
      \-vma18\   : in  std_logic;
      \-vmo19\   : out std_logic;
      \-vma19\   : in  std_logic;
      \-vmo12\   : out std_logic;
      \-vma12\   : in  std_logic;
      \-vmo13\   : out std_logic;
      \-vma13\   : in  std_logic;
      \-vmo14\   : out std_logic;
      \-vma14\   : in  std_logic;
      \-vmo15\   : out std_logic;
      \-vma15\   : in  std_logic;
      vmoparm    : out std_logic;
      vmopar     : out std_logic;
      vm1pari    : in  std_logic;
      \-vmap4\   : in  std_logic;
      \-vmap3\   : in  std_logic;
      \-vmap2\   : in  std_logic;
      \-vmap1\   : in  std_logic;
      \-vmap0\   : in  std_logic;
      \-vmo5\    : in  std_logic;
      \-vmo6\    : in  std_logic;
      \-vmo7\    : in  std_logic;
      \-vmo8\    : in  std_logic;
      \-vmo9\    : in  std_logic;
      \-vmo10\   : in  std_logic;
      \-vmo11\   : in  std_logic;
      vmoparl    : out std_logic;
      \-vmo0\    : in  std_logic;
      \-vmo1\    : in  std_logic;
      \-vmo2\    : in  std_logic;
      \-vmo3\    : in  std_logic;
      \-vmo4\    : in  std_logic;
      vmoparodd  : out std_logic;
      vmoparck   : out std_logic
      );
  end component;

  component cadr_vmemdr is
    port (
      \-mapdrive\ : out std_logic;
      \-pfw\      : in  std_logic;
      mf24        : out std_logic;
      \-pfr\      : in  std_logic;
      mf25        : out std_logic;
      mf26        : out std_logic;
      \-vmap4\    : in  std_logic;
      mf27        : out std_logic;
      \-vmap3\    : in  std_logic;
      mf28        : out std_logic;
      \-vmap2\    : in  std_logic;
      mf29        : out std_logic;
      \-vmap1\    : in  std_logic;
      mf30        : out std_logic;
      \-vmap0\    : in  std_logic;
      mf31        : out std_logic;
      \-vmo15\    : in  std_logic;
      mf8         : out std_logic;
      \-vmo14\    : in  std_logic;
      mf9         : out std_logic;
      \-vmo13\    : in  std_logic;
      mf10        : out std_logic;
      \-vmo12\    : in  std_logic;
      mf11        : out std_logic;
      \-vmo11\    : in  std_logic;
      mf12        : out std_logic;
      \-vmo10\    : in  std_logic;
      mf13        : out std_logic;
      \-vmo9\     : in  std_logic;
      mf14        : out std_logic;
      \-vmo8\     : in  std_logic;
      mf15        : out std_logic;
      \-vmo23\    : in  std_logic;
      mf16        : out std_logic;
      \-vmo22\    : in  std_logic;
      mf17        : out std_logic;
      \-vmo21\    : in  std_logic;
      mf18        : out std_logic;
      \-vmo20\    : in  std_logic;
      mf19        : out std_logic;
      \-vmo19\    : in  std_logic;
      mf20        : out std_logic;
      \-vmo18\    : in  std_logic;
      mf21        : out std_logic;
      \-vmo17\    : in  std_logic;
      mf22        : out std_logic;
      \-vmo16\    : in  std_logic;
      mf23        : out std_logic;
      tse1a       : in  std_logic;
      srcmap      : out std_logic;
      \-vmo7\     : in  std_logic;
      mf0         : out std_logic;
      \-vmo6\     : in  std_logic;
      mf1         : out std_logic;
      \-vmo5\     : in  std_logic;
      mf2         : out std_logic;
      \-vmo4\     : in  std_logic;
      mf3         : out std_logic;
      \-vmo3\     : in  std_logic;
      mf4         : out std_logic;
      \-vmo2\     : in  std_logic;
      mf5         : out std_logic;
      \-vmo1\     : in  std_logic;
      mf6         : out std_logic;
      \-vmo0\     : in  std_logic;
      mf7         : out std_logic;
      \-lvmo23\   : out std_logic;
      \-lvmo22\   : out std_logic;
      \-pma21\    : out std_logic;
      \-pma20\    : out std_logic;
      memstart    : in  std_logic;
      \-pma19\    : out std_logic;
      \-pma18\    : out std_logic;
      \-pma17\    : out std_logic;
      \-pma16\    : out std_logic;
      \-pma15\    : out std_logic;
      \-pma14\    : out std_logic;
      \-pma13\    : out std_logic;
      \-pma12\    : out std_logic;
      \-pma11\    : out std_logic;
      \-pma10\    : out std_logic;
      \-pma9\     : out std_logic;
      \-pma8\     : out std_logic;
      \-vma6\     : in  std_logic;
      \-vma5\     : in  std_logic;
      \-vma4\     : in  std_logic;
      \-vma3\     : in  std_logic;
      \-vma2\     : in  std_logic;
      \-vma1\     : in  std_logic;
      \-vma0\     : in  std_logic;
      \-vma7\     : in  std_logic;
      \-adrpar\   : out std_logic;
      \-srcmap\   : in  std_logic
      );
  end component;

end package;

