library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_q is
  port (
    hi7      : in  std_logic;
    q23      : out std_logic;
    alu24    : in  std_logic;
    alu25    : in  std_logic;
    alu26    : in  std_logic;
    alu27    : in  std_logic;
    q28      : out std_logic;
    qs0      : in  std_logic;
    qs1      : in  std_logic;
    clk2b    : in  std_logic;
    q27      : out std_logic;
    q26      : out std_logic;
    q25      : out std_logic;
    q24      : out std_logic;
    alu28    : in  std_logic;
    alu29    : in  std_logic;
    alu30    : in  std_logic;
    alu31    : in  std_logic;
    alu0     : in  std_logic;
    q31      : out std_logic;
    q30      : out std_logic;
    q29      : out std_logic;
    q15      : out std_logic;
    alu16    : in  std_logic;
    alu17    : in  std_logic;
    alu18    : in  std_logic;
    alu19    : in  std_logic;
    q20      : out std_logic;
    q19      : out std_logic;
    q18      : out std_logic;
    q17      : out std_logic;
    q16      : out std_logic;
    alu20    : in  std_logic;
    alu21    : in  std_logic;
    alu22    : in  std_logic;
    alu23    : in  std_logic;
    q22      : out std_logic;
    q21      : out std_logic;
    q7       : out std_logic;
    alu8     : in  std_logic;
    alu9     : in  std_logic;
    alu10    : in  std_logic;
    alu11    : in  std_logic;
    q12      : out std_logic;
    q11      : out std_logic;
    q10      : out std_logic;
    q9       : out std_logic;
    q8       : out std_logic;
    alu12    : in  std_logic;
    alu13    : in  std_logic;
    alu14    : in  std_logic;
    alu15    : in  std_logic;
    q14      : out std_logic;
    q13      : out std_logic;
    \-alu31\ : in  std_logic;
    alu1     : in  std_logic;
    alu2     : in  std_logic;
    alu3     : in  std_logic;
    q4       : out std_logic;
    q3       : out std_logic;
    q2       : out std_logic;
    q1       : out std_logic;
    q0       : out std_logic;
    alu4     : in  std_logic;
    alu5     : in  std_logic;
    alu6     : in  std_logic;
    alu7     : in  std_logic;
    q6       : out std_logic;
    q5       : out std_logic);
end;

architecture ttl of cadr4_q is
begin
  q_2c07 : sn74s194 port map(clr_n => hi7, sir => q23, i0 => alu24, i1 => alu25, i2 => alu26, i3 => alu27, sil => q28, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q27, q2 => q26, q1 => q25, q0 => q24);
  q_2c08 : sn74s194 port map(clr_n => hi7, sir => q27, i0 => alu28, i1 => alu29, i2 => alu30, i3 => alu31, sil => alu0, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q31, q2 => q30, q1 => q29, q0 => q28);
  q_2c12 : sn74s194 port map(clr_n => hi7, sir => q15, i0 => alu16, i1 => alu17, i2 => alu18, i3 => alu19, sil => q20, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q19, q2 => q18, q1 => q17, q0 => q16);
  q_2c13 : sn74s194 port map(clr_n => hi7, sir => q19, i0 => alu20, i1 => alu21, i2 => alu22, i3 => alu23, sil => q24, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q23, q2 => q22, q1 => q21, q0 => q20);
  q_2c22 : sn74s194 port map(clr_n => hi7, sir => q7, i0 => alu8, i1 => alu9, i2 => alu10, i3 => alu11, sil => q12, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q11, q2 => q10, q1 => q9, q0 => q8);
  q_2c23 : sn74s194 port map(clr_n => hi7, sir => q11, i0 => alu12, i1 => alu13, i2 => alu14, i3 => alu15, sil => q16, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q15, q2 => q14, q1 => q13, q0 => q12);
  q_2c27 : sn74s194 port map(clr_n => hi7, sir => \-alu31\, i0 => alu0, i1 => alu1, i2 => alu2, i3 => alu3, sil => q4, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q3, q2 => q2, q1 => q1, q0 => q0);
  q_2c28 : sn74s194 port map(clr_n => hi7, sir => q3, i0 => alu4, i1 => alu5, i2 => alu6, i3 => alu7, sil => q8, s0 => qs0, s1 => qs1, clk => clk2b, q3 => q7, q2 => q6, q1 => q5, q0 => q4);
end architecture;
