library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_ictl is
  port (
    ramdisable      : out std_logic;
    hi1             : in  std_logic;
    \-iwriteda\     : out std_logic;
    \-promdisabled\ : out std_logic;
    idebug          : in  std_logic;
    iwriteda        : out std_logic;
    promdisabled    : in  std_logic;
    \-wp5\          : in  std_logic;
    wp5d            : out std_logic;
    wp5c            : out std_logic;
    wp5b            : out std_logic;
    wp5a            : out std_logic;
    pc0             : in  std_logic;
    \-pcb0\         : out std_logic;
    pc1             : in  std_logic;
    \-pcb1\         : out std_logic;
    pc2             : in  std_logic;
    \-pcb2\         : out std_logic;
    \-pcb3\         : out std_logic;
    pc3             : in  std_logic;
    \-pcb4\         : out std_logic;
    pc4             : in  std_logic;
    \-pcb5\         : out std_logic;
    pc5             : in  std_logic;
    \-iwea\         : out std_logic;
    \-iweb\         : out std_logic;
    \-iwei\         : out std_logic;
    \-iwej\         : out std_logic;
    pc13            : in  std_logic;
    \-pc13b\        : out std_logic;
    pc12            : in  std_logic;
    \-pc12b\        : out std_logic;
    \-iwrited\      : in  std_logic;
    iwritedd        : out std_logic;
    iwritedc        : out std_logic;
    iwritedb        : out std_logic;
    pc6             : in  std_logic;
    \-pcb6\         : out std_logic;
    pc7             : in  std_logic;
    \-pcb7\         : out std_logic;
    pc8             : in  std_logic;
    \-pcb8\         : out std_logic;
    \-pcb9\         : out std_logic;
    pc9             : in  std_logic;
    \-pcb10\        : out std_logic;
    pc10            : in  std_logic;
    \-pcb11\        : out std_logic;
    pc11            : in  std_logic;
    \-ice3a\        : out std_logic;
    \-ice2a\        : out std_logic;
    \-ice1a\        : out std_logic;
    \-ice0a\        : out std_logic;
    \-ice0b\        : out std_logic;
    \-ice1b\        : out std_logic;
    \-ice2b\        : out std_logic;
    \-ice3b\        : out std_logic;
    \-iwec\         : out std_logic;
    \-iwed\         : out std_logic;
    \-iwek\         : out std_logic;
    \-iwel\         : out std_logic;
    \-pcc0\         : out std_logic;
    \-pcc1\         : out std_logic;
    \-pcc2\         : out std_logic;
    \-pcc3\         : out std_logic;
    \-pcc4\         : out std_logic;
    \-pcc5\         : out std_logic;
    \-pcc6\         : out std_logic;
    \-pcc7\         : out std_logic;
    \-pcc8\         : out std_logic;
    \-pcc9\         : out std_logic;
    \-pcc10\        : out std_logic;
    \-pcc11\        : out std_logic;
    \-iwee\         : out std_logic;
    \-iwef\         : out std_logic;
    \-iwem\         : out std_logic;
    \-iwen\         : out std_logic;
    \-ice3c\        : out std_logic;
    \-ice2c\        : out std_logic;
    \-ice1c\        : out std_logic;
    \-ice0c\        : out std_logic;
    \-ice0d\        : out std_logic;
    \-ice1d\        : out std_logic;
    \-ice2d\        : out std_logic;
    \-ice3d\        : out std_logic;
    \-iweg\         : out std_logic;
    \-iweh\         : out std_logic;
    \-iweo\         : out std_logic;
    \-iwep\         : out std_logic);
end;

architecture ttl of cadr4_ictl is
begin
  ictl_1a15 : dm9s42_1 port map(out2 => ramdisable, g2d2 => hi1, g2c2 => hi1, g2b2 => \-iwriteda\, g2a2 => \-promdisabled\, g1b2 => hi1, g1a2 => idebug, g1a1 => '0', g1b1 => '0', g2a1 => '0', g2b1 => '0', g2c1 => '0', g2d1 => '0');
  ictl_1c16 : sn74s04 port map(g1a   => iwriteda, g1q_n => \-iwriteda\, g2a => promdisabled, g2q_n => \-promdisabled\, g3a => \-wp5\, g3q_n => wp5d, g4q_n => wp5c, g4a => \-wp5\, g5q_n => wp5b, g5a => \-wp5\, g6q_n => wp5a, g6a => \-wp5\);
  ictl_1c21 : sn74s04 port map(g1a   => pc0, g1q_n => \-pcb0\, g2a => pc1, g2q_n => \-pcb1\, g3a => pc2, g3q_n => \-pcb2\, g4q_n => \-pcb3\, g4a => pc3, g5q_n => \-pcb4\, g5a => pc4, g6q_n => \-pcb5\, g6a => pc5);
  ictl_1c26 : sn74s37 port map(g1a   => wp5a, g1b => iwriteda, g1y => \-iwea\, g2a => wp5a, g2b => iwriteda, g2y => \-iweb\, g3y => \-iwei\, g3a => iwriteda, g3b => wp5a, g4y => \-iwej\, g4a => iwriteda, g4b => wp5a);
  ictl_1d20 : sn74s04 port map(g1a   => pc13, g1q_n => \-pc13b\, g2a => pc12, g2q_n => \-pc12b\, g3a => \-iwrited\, g3q_n => iwritedd, g4q_n => iwritedc, g4a => \-iwrited\, g5q_n => iwritedb, g5a => \-iwrited\, g6q_n => iwriteda, g6a => \-iwrited\);
  ictl_1d25 : sn74s04 port map(g1a   => pc6, g1q_n => \-pcb6\, g2a => pc7, g2q_n => \-pcb7\, g3a => pc8, g3q_n => \-pcb8\, g4q_n => \-pcb9\, g4a => pc9, g5q_n => \-pcb10\, g5a => pc10, g6q_n => \-pcb11\, g6a => pc11);
  ictl_1d30 : sn74s139 port map(g1   => ramdisable, a1 => \-pc12b\, b1 => \-pc13b\, g1y0 => \-ice3a\, g1y1 => \-ice2a\, g1y2 => \-ice1a\, g1y3 => \-ice0a\, g2y3 => \-ice0b\, g2y2 => \-ice1b\, g2y1 => \-ice2b\, g2y0 => \-ice3b\, b2 => \-pc13b\, a2 => \-pc12b\, g2 => ramdisable);
  ictl_2c01 : sn74s37 port map(g1a   => wp5b, g1b => iwritedb, g1y => \-iwec\, g2a => wp5b, g2b => iwritedb, g2y => \-iwed\, g3y => \-iwek\, g3a => iwritedb, g3b => wp5b, g4y => \-iwel\, g4a => iwritedb, g4b => wp5b);
  ictl_2c06 : sn74s04 port map(g1a   => pc0, g1q_n => \-pcc0\, g2a => pc1, g2q_n => \-pcc1\, g3a => pc2, g3q_n => \-pcc2\, g4q_n => \-pcc3\, g4a => pc3, g5q_n => \-pcc4\, g5a => pc4, g6q_n => \-pcc5\, g6a => pc5);
  ictl_2d10 : sn74s04 port map(g1a   => pc6, g1q_n => \-pcc6\, g2a => pc7, g2q_n => \-pcc7\, g3a => pc8, g3q_n => \-pcc8\, g4q_n => \-pcc9\, g4a => pc9, g5q_n => \-pcc10\, g5a => pc10, g6q_n => \-pcc11\, g6a => pc11);
  ictl_2d15 : sn74s37 port map(g1a   => wp5c, g1b => iwritedc, g1y => \-iwee\, g2a => wp5c, g2b => iwritedc, g2y => \-iwef\, g3y => \-iwem\, g3a => iwritedc, g3b => wp5c, g4y => \-iwen\, g4a => iwritedc, g4b => wp5c);
  ictl_2d25 : sn74s139 port map(g1   => ramdisable, a1 => \-pc12b\, b1 => \-pc13b\, g1y0 => \-ice3c\, g1y1 => \-ice2c\, g1y2 => \-ice1c\, g1y3 => \-ice0c\, g2y3 => \-ice0d\, g2y2 => \-ice1d\, g2y1 => \-ice2d\, g2y0 => \-ice3d\, b2 => \-pc13b\, a2 => \-pc12b\, g2 => ramdisable);
  ictl_2d30 : sn74s37 port map(g1a   => wp5d, g1b => iwritedd, g1y => \-iweg\, g2a => wp5d, g2b => iwritedd, g2y => \-iweh\, g3y => \-iweo\, g3a => iwritedd, g3b => wp5d, g4y => \-iwep\, g4a => iwritedd, g4b => wp5d);
end architecture;
