-- CADR1_LMADR
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_lmadr is
  port (
    \-adr0\ : inout std_logic;
    \-adr1\ : inout std_logic;
    \-adr10\ : inout std_logic;
    \-adr11\ : inout std_logic;
    \-adr12\ : inout std_logic;
    \-adr13\ : inout std_logic;
    \-adr14\ : inout std_logic;
    \-adr15\ : inout std_logic;
    \-adr16\ : inout std_logic;
    \-adr17\ : inout std_logic;
    \-adr18\ : inout std_logic;
    \-adr19\ : inout std_logic;
    \-adr2\ : inout std_logic;
    \-adr3\ : inout std_logic;
    \-adr4\ : inout std_logic;
    \-adr5\ : inout std_logic;
    \-adr6\ : inout std_logic;
    \-adr7\ : inout std_logic;
    \-adr8\ : inout std_logic;
    \-adr9\ : inout std_logic;
    \-lmadr_ub\ : inout std_logic;
    \-lmadr_xbus\ : inout std_logic;
    uao1 : inout std_logic;
    uao10 : inout std_logic;
    uao11 : inout std_logic;
    uao12 : inout std_logic;
    uao13 : inout std_logic;
    uao14 : inout std_logic;
    uao15 : inout std_logic;
    uao16 : inout std_logic;
    uao17 : inout std_logic;
    uao2 : inout std_logic;
    uao3 : inout std_logic;
    uao4 : inout std_logic;
    uao5 : inout std_logic;
    uao6 : inout std_logic;
    uao7 : inout std_logic;
    uao8 : inout std_logic;
    uao9 : inout std_logic;
    xao0 : inout std_logic;
    xao1 : inout std_logic;
    xao10 : inout std_logic;
    xao11 : inout std_logic;
    xao12 : inout std_logic;
    xao13 : inout std_logic;
    xao14 : inout std_logic;
    xao15 : inout std_logic;
    xao16 : inout std_logic;
    xao17 : inout std_logic;
    xao18 : inout std_logic;
    xao19 : inout std_logic;
    xao2 : inout std_logic;
    xao3 : inout std_logic;
    xao4 : inout std_logic;
    xao5 : inout std_logic;
    xao6 : inout std_logic;
    xao7 : inout std_logic;
    xao8 : inout std_logic;
    xao9 : inout std_logic
  );
end entity;
