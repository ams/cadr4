library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_mf is
  port (
    tse1a      : in  std_logic;
    mfenb      : out std_logic;
    \-mfdrive\ : out std_logic;
    mf23       : in  std_logic;
    m16        : out std_logic;
    mf22       : in  std_logic;
    m17        : out std_logic;
    mf21       : in  std_logic;
    m18        : out std_logic;
    mf20       : in  std_logic;
    m19        : out std_logic;
    mf19       : in  std_logic;
    m20        : out std_logic;
    mf18       : in  std_logic;
    m21        : out std_logic;
    mf17       : in  std_logic;
    m22        : out std_logic;
    mf16       : in  std_logic;
    m23        : out std_logic;
    mfdrive    : out std_logic;
    mf15       : in  std_logic;
    m8         : out std_logic;
    mf14       : in  std_logic;
    m9         : out std_logic;
    mf13       : in  std_logic;
    m10        : out std_logic;
    mf12       : in  std_logic;
    m11        : out std_logic;
    mf11       : in  std_logic;
    m12        : out std_logic;
    mf10       : in  std_logic;
    m13        : out std_logic;
    mf9        : in  std_logic;
    m14        : out std_logic;
    mf8        : in  std_logic;
    m15        : out std_logic;
    mf7        : in  std_logic;
    m0         : out std_logic;
    mf6        : in  std_logic;
    m1         : out std_logic;
    mf5        : in  std_logic;
    m2         : out std_logic;
    mf4        : in  std_logic;
    m3         : out std_logic;
    mf3        : in  std_logic;
    m4         : out std_logic;
    mf2        : in  std_logic;
    m5         : out std_logic;
    mf1        : in  std_logic;
    m6         : out std_logic;
    mf0        : in  std_logic;
    m7         : out std_logic;
    mf31       : in  std_logic;
    m24        : out std_logic;
    mf30       : in  std_logic;
    m25        : out std_logic;
    mf29       : in  std_logic;
    m26        : out std_logic;
    mf28       : in  std_logic;
    m27        : out std_logic;
    mf27       : in  std_logic;
    m28        : out std_logic;
    mf26       : in  std_logic;
    m29        : out std_logic;
    mf25       : in  std_logic;
    m30        : out std_logic;
    mf24       : in  std_logic;
    m31        : out std_logic;
    pdlenb     : in  std_logic;
    spcenb     : in  std_logic;
    \-srcm\    : out std_logic;
    \-ir31\    : in  std_logic;
    \-mpass\   : in  std_logic);
end;

architecture ttl of cadr_mf is
  signal internal22 : std_logic;
begin
  mf_1a18 : sn74s00 port map(g1b     => tse1a, g1a => mfenb, g1q_n => \-mfdrive\, g2b => '0', g2a => '0', g3b => '0', g3a => '0', g4a => '0', g4b => '0');
  mf_1a21 : sn74s241 port map(aenb_n => \-mfdrive\, ain0 => mf23, bout3 => m16, ain1 => mf22, bout2 => m17, ain2 => mf21, bout1 => m18, ain3 => mf20, bout0 => m19, bin0 => mf19, aout3 => m20, bin1 => mf18, aout2 => m21, bin2 => mf17, aout1 => m22, bin3 => mf16, aout0 => m23, benb => mfdrive);
  mf_1a23 : sn74s241 port map(aenb_n => \-mfdrive\, ain0 => mf15, bout3 => m8, ain1 => mf14, bout2 => m9, ain2 => mf13, bout1 => m10, ain3 => mf12, bout0 => m11, bin0 => mf11, aout3 => m12, bin1 => mf10, aout2 => m13, bin2 => mf9, aout1 => m14, bin3 => mf8, aout0 => m15, benb => mfdrive);
  mf_1a25 : sn74s241 port map(aenb_n => \-mfdrive\, ain0 => mf7, bout3 => m0, ain1 => mf6, bout2 => m1, ain2 => mf5, bout1 => m2, ain3 => mf4, bout0 => m3, bin0 => mf3, aout3 => m4, bin1 => mf2, aout2 => m5, bin2 => mf1, aout1 => m6, bin3 => mf0, aout0 => m7, benb => mfdrive);
  mf_1b24 : sn74s241 port map(aenb_n => \-mfdrive\, ain0 => mf31, bout3 => m24, ain1 => mf30, bout2 => m25, ain2 => mf29, bout1 => m26, ain3 => mf28, bout0 => m27, bin0 => mf27, aout3 => m28, bin1 => mf26, aout2 => m29, bin2 => mf25, aout1 => m30, bin3 => mf24, aout0 => m31, benb => mfdrive);
  mf_2a04 : sn74s08 port map(g2b     => tse1a, g2a => mfenb, g2q => mfdrive, g1b => '0', g1a => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  mf_3f14 : sn74s02 port map(g3b     => pdlenb, g3a => spcenb, g3q_n => internal22, g1a => '0', g1b => '0', g2a => '0', g2b => '0', g4b => '0', g4a => '0');
  mf_4d06 : sn74s08 port map(g4q     => mfenb, g4a => internal22, g4b => \-srcm\, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3a => '0', g3b => '0');
  mf_4d08 : sn74s00 port map(g4q_n   => \-srcm\, g4a => \-ir31\, g4b => \-mpass\, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3b => '0', g3a => '0');
end architecture;
