library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_l is
  port (
    gnd        : in  std_logic;
    l7         : out std_logic;
    ob7        : in  std_logic;
    ob6        : in  std_logic;
    l6         : out std_logic;
    l5         : out std_logic;
    ob5        : in  std_logic;
    ob4        : in  std_logic;
    l4         : out std_logic;
    clk3f      : in  std_logic;
    l3         : out std_logic;
    ob3        : in  std_logic;
    ob2        : in  std_logic;
    l2         : out std_logic;
    l1         : out std_logic;
    ob1        : in  std_logic;
    ob0        : in  std_logic;
    l0         : out std_logic;
    l15        : out std_logic;
    ob15       : in  std_logic;
    ob14       : in  std_logic;
    l14        : out std_logic;
    l13        : out std_logic;
    ob13       : in  std_logic;
    ob12       : in  std_logic;
    l12        : out std_logic;
    l11        : out std_logic;
    ob11       : in  std_logic;
    ob10       : in  std_logic;
    l10        : out std_logic;
    l9         : out std_logic;
    ob9        : in  std_logic;
    ob8        : in  std_logic;
    l8         : out std_logic;
    l23        : out std_logic;
    ob23       : in  std_logic;
    ob22       : in  std_logic;
    l22        : out std_logic;
    l21        : out std_logic;
    ob21       : in  std_logic;
    ob20       : in  std_logic;
    l20        : out std_logic;
    l19        : out std_logic;
    ob19       : in  std_logic;
    ob18       : in  std_logic;
    l18        : out std_logic;
    l17        : out std_logic;
    ob17       : in  std_logic;
    ob16       : in  std_logic;
    l16        : out std_logic;
    l31        : out std_logic;
    ob31       : in  std_logic;
    ob30       : in  std_logic;
    l30        : out std_logic;
    l29        : out std_logic;
    ob29       : in  std_logic;
    ob28       : in  std_logic;
    l28        : out std_logic;
    l27        : out std_logic;
    ob27       : in  std_logic;
    ob26       : in  std_logic;
    l26        : out std_logic;
    l25        : out std_logic;
    ob25       : in  std_logic;
    ob24       : in  std_logic;
    l24        : out std_logic;
    lparl      : out std_logic;
    nc369      : out std_logic;
    nc370      : out std_logic;
    \-lparm\   : out std_logic;
    lparity    : out std_logic;
    \-lparity\ : out std_logic);
end;

architecture ttl of cadr4_l is
begin
  l_3c26 : sn74s374 port map(oenb_n => gnd, o0 => l7, i0 => ob7, i1 => ob6, o1 => l6, o2 => l5, i2 => ob5, i3 => ob4, o3 => l4, clk => clk3f, o4 => l3, i4 => ob3, i5 => ob2, o5 => l2, o6 => l1, i6 => ob1, i7 => ob0, o7 => l0);
  l_3c27 : sn74s374 port map(oenb_n => gnd, o0 => l15, i0 => ob15, i1 => ob14, o1 => l14, o2 => l13, i2 => ob13, i3 => ob12, o3 => l12, clk => clk3f, o4 => l11, i4 => ob11, i5 => ob10, o5 => l10, o6 => l9, i6 => ob9, i7 => ob8, o7 => l8);
  l_3c28 : sn74s374 port map(oenb_n => gnd, o0 => l23, i0 => ob23, i1 => ob22, o1 => l22, o2 => l21, i2 => ob21, i3 => ob20, o3 => l20, clk => clk3f, o4 => l19, i4 => ob19, i5 => ob18, o5 => l18, o6 => l17, i6 => ob17, i7 => ob16, o7 => l16);
  l_3c29 : sn74s374 port map(oenb_n => gnd, o0 => l31, i0 => ob31, i1 => ob30, o1 => l30, o2 => l29, i2 => ob29, i3 => ob28, o3 => l28, clk => clk3f, o4 => l27, i4 => ob27, i5 => ob26, o5 => l26, o6 => l25, i6 => ob25, i7 => ob24, o7 => l24);
  l_4c03 : am93s48 port map(i6      => l5, i5 => l6, i4 => l7, i3 => l8, i2 => l9, i1 => l10, i0 => l11, po => lparl, pe => nc369, i11 => l0, i10 => l1, i9 => l2, i8 => l3, i7 => l4);
  l_4c08 : am93s48 port map(i6      => l17, i5 => l18, i4 => l19, i3 => l20, i2 => l21, i1 => l22, i0 => l23, po => nc370, pe => \-lparm\, i11 => l12, i10 => l13, i9 => l14, i8 => l15, i7 => l16);
  l_4c09 : am93s48 port map(i6      => l25, i5 => l26, i4 => l27, i3 => l28, i2 => l29, i1 => l30, i0 => l31, po => lparity, pe => \-lparity\, i11 => lparl, i10 => \-lparm\, i9 => gnd, i8 => gnd, i7 => l24);
end architecture;
