library ieee;
use ieee.std_logic_1164.all;

-- Dec 14 18:19:44 1980

package cadr_book is

  component actl is
    port ();
  end component;

  component alatch is
    port ();
  end component;

  component alu0 is
    port ();
  end component;

  component alu1 is
    port ();
  end component;

  component aluc4 is
    port ();
  end component;

  component amem0 is
    port ();
  end component;

  component amem1 is
    port ();
  end component;

  component apar is
    port ();
  end component;

  component bcpins is
    port ();
  end component;

  component bcterm is
    port ();
  end component;

  component caps is
    port ();
  end component;

  component clockd is
    port ();
  end component;

  component contrl is
    port ();
  end component;

  component cpins is
    port ();
  end component;

  component dram0 is
    port ();
  end component;

  component dram1 is
    port ();
  end component;

  component dram2 is
    port ();
  end component;

  component dspctl is
    port ();
  end component;

  component flag is
    port ();
  end component;

  component ior is
    port ();
  end component;

  component ipar is
    port ();
  end component;

  component ireg is
    port ();
  end component;

  component iwr is
    port ();
  end component;

  component l is
    port ();
  end component;

  component lc is
    port ();
  end component;

  component lcc is
    port ();
  end component;

  component lpc is
    port ();
  end component;

  component mctl is
    port ();
  end component;

  component md is
    port ();
  end component;

  component mds is
    port ();
  end component;

  component mf is
    port ();
  end component;

  component mlatch is
    port ();
  end component;

  component mmem is
    port ();
  end component;

  component mo0 is
    port ();
  end component;

  component mo1 is
    port ();
  end component;

  component mskg4 is
    port ();
  end component;

  component npc is
    port ();
  end component;

  component opcd is
    port ();
  end component;

  component pdl0 is
    port ();
  end component;

  component pdl1 is
    port ();
  end component;

  component pdlctl is
    port ();
  end component;

  component pdlptr is
    port ();
  end component;

  component platch is
    port ();
  end component;

  component q is
    port ();
  end component;

  component qctl is
    port ();
  end component;

  component shift0 is
    port ();
  end component;

  component shift1 is
    port ();
  end component;

  component smctl is
    port ();
  end component;

  component source is
    port ();
  end component;

  component spc is
    port ();
  end component;

  component spclch is
    port ();
  end component;

  component spcpar is
    port ();
  end component;

  component spcw is
    port ();
  end component;

  component spy1 is
    port ();
  end component;

  component spy2 is
    port ();
  end component;

  component trap is
    port ();
  end component;

  component vctl1 is
    port ();
  end component;

  component vctl2 is
    port ();
  end component;

  component vma is
    port ();
  end component;

  component vmas is
    port ();
  end component;

  component vmem0 is
    port ();
  end component;

  component vmem1 is
    port ();
  end component;

  component vmem2 is
    port ();
  end component;

  component vmemdr is
    port ();
  end component;

end package;
