library ieee;
use ieee.std_logic_1164.all;

entity cadr_pctl is
  port (
    \-promenable\   : out std_logic;
    i46             : out std_logic;
    hi2             : in  std_logic;
    pc0             : in  std_logic;
    \-prompc0\      : out std_logic;
    pc1             : in  std_logic;
    \-prompc1\      : out std_logic;
    pc2             : in  std_logic;
    \-prompc2\      : out std_logic;
    \-prompc3\      : out std_logic;
    pc3             : in  std_logic;
    \-prompc4\      : out std_logic;
    pc4             : in  std_logic;
    pc9             : in  std_logic;
    \-promce0\      : out std_logic;
    \-prompc9\      : out std_logic;
    \-promce1\      : out std_logic;
    \bottom.1k\     : out std_logic;
    \-idebug\       : in  std_logic;
    \-promdisabled\ : in  std_logic;
    \-iwriteda\     : in  std_logic;
    pc13            : in  std_logic;
    pc11            : in  std_logic;
    pc10            : in  std_logic;
    pc5             : in  std_logic;
    \-prompc5\      : out std_logic;
    pc6             : in  std_logic;
    \-prompc6\      : out std_logic;
    pc7             : in  std_logic;
    \-prompc7\      : out std_logic;
    \-prompc8\      : out std_logic;
    pc8             : in  std_logic;
    \-ape\          : in  std_logic;
    \-pdlpe\        : in  std_logic;
    \-spe\          : in  std_logic;
    \-mpe\          : in  std_logic;
    tilt1           : out std_logic;
    tilt0           : out std_logic;
    \-mempe\        : in  std_logic;
    \-v1pe\         : in  std_logic;
    \-v0pe\         : in  std_logic;
    promenable      : out std_logic;
    dpe             : out std_logic;
    \-dpe\          : in  std_logic;
    ipe             : out std_logic;
    \-ipe\          : in  std_logic;
    pc12            : in  std_logic
    );
end;
