library ieee;
use ieee.std_logic_1164.all;

entity cadr_spc is
  port (
    \-swpa\   : in  std_logic;
    spcw14    : in  std_logic;
    spcptr4   : out std_logic;
    spco14    : out std_logic;
    spco15    : out std_logic;
    spcptr3   : out std_logic;
    spcptr2   : out std_logic;
    spcptr1   : out std_logic;
    spcptr0   : out std_logic;
    spcw15    : in  std_logic;
    spcw12    : in  std_logic;
    spco12    : out std_logic;
    spco13    : out std_logic;
    spcw13    : in  std_logic;
    spcw10    : in  std_logic;
    spco10    : out std_logic;
    spco11    : out std_logic;
    spcw11    : in  std_logic;
    spcopar   : out std_logic;
    spco18    : out std_logic;
    spco17    : out std_logic;
    spco16    : out std_logic;
    \-swpb\   : in  std_logic;
    spcw4     : in  std_logic;
    spco4     : out std_logic;
    spco5     : out std_logic;
    spcw5     : in  std_logic;
    spcw2     : in  std_logic;
    spco2     : out std_logic;
    spco3     : out std_logic;
    spcw3     : in  std_logic;
    spcw0     : in  std_logic;
    spco0     : out std_logic;
    spco1     : out std_logic;
    spcw1     : in  std_logic;
    spco9     : out std_logic;
    spco8     : out std_logic;
    spco7     : out std_logic;
    spco6     : out std_logic;
    spush     : in  std_logic;
    clk4f     : in  std_logic;
    \-spcnt\  : in  std_logic;
    \-spccry\ : out std_logic;
    spcw18    : in  std_logic;
    spcwpar   : in  std_logic;
    spcw16    : in  std_logic;
    spcw17    : in  std_logic;
    spcw8     : in  std_logic;
    spcw9     : in  std_logic;
    spcw6     : in  std_logic;
    spcw7     : in  std_logic
    );
end;
