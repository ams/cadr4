-- D Flip-Flop

library ieee;
use ieee.std_logic_1164.all;

entity ff_d is
  port (
    clk    : in  std_logic := 'H';
    d      : in  std_logic := 'H';
    enb_n  : in  std_logic := '0';
    q, q_n : out std_logic
    );
end;

architecture ttl of ff_d is
  signal q_int : std_logic;
begin

  q <= q_int;
  -- Proper complement handling for unknown states
  q_n <= '0' when q_int = '1' else
         '1' when q_int = '0' else
         'X';  -- Unknown complement for X, U, Z, W states

  process (clk)
  begin
    if to_x01(enb_n) = '0' then
      -- Handle metavalue clock transitions
      if clk'event then
        if is_x(clk) or is_x(clk'last_value) then
          -- Clock transition involving metavalue - output becomes unknown
          q_int <= 'X';
        elsif clk = '1' and clk'last_value = '0' then
          -- Valid rising edge
          q_int <= d;
        end if;
      end if;
    end if;
  end process;

end;
