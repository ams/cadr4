library ieee;
use ieee.std_logic_1164.all;

entity cadr_spc is
  port (
    \-spcnt\        : in     std_logic;
    \-swpa\         : in     std_logic;
    \-swpb\         : in     std_logic;
    clk4f           : in     std_logic;
    spcw0           : in     std_logic;
    spcw1           : in     std_logic;
    spcw10          : in     std_logic;
    spcw11          : in     std_logic;
    spcw12          : in     std_logic;
    spcw13          : in     std_logic;
    spcw14          : in     std_logic;
    spcw15          : in     std_logic;
    spcw16          : in     std_logic;
    spcw17          : in     std_logic;
    spcw18          : in     std_logic;
    spcw2           : in     std_logic;
    spcw3           : in     std_logic;
    spcw4           : in     std_logic;
    spcw5           : in     std_logic;
    spcw6           : in     std_logic;
    spcw7           : in     std_logic;
    spcw8           : in     std_logic;
    spcw9           : in     std_logic;
    spcwpar         : in     std_logic;
    spush           : in     std_logic;
    hi1             : inout  std_logic;
    hi10            : inout  std_logic;
    hi11            : inout  std_logic;
    hi12            : inout  std_logic;
    hi2             : inout  std_logic;
    hi3             : inout  std_logic;
    hi4             : inout  std_logic;
    hi5             : inout  std_logic;
    hi6             : inout  std_logic;
    hi7             : inout  std_logic;
    hi8             : inout  std_logic;
    hi9             : inout  std_logic;
    spco0           : inout  std_logic;
    spco1           : inout  std_logic;
    spco10          : inout  std_logic;
    spco11          : inout  std_logic;
    spco12          : inout  std_logic;
    spco13          : inout  std_logic;
    spco14          : inout  std_logic;
    spco15          : inout  std_logic;
    spco16          : inout  std_logic;
    spco17          : inout  std_logic;
    spco18          : inout  std_logic;
    spco2           : inout  std_logic;
    spco3           : inout  std_logic;
    spco4           : inout  std_logic;
    spco5           : inout  std_logic;
    spco6           : inout  std_logic;
    spco7           : inout  std_logic;
    spco8           : inout  std_logic;
    spco9           : inout  std_logic;
    spcopar         : inout  std_logic;
    \-spccry\       : out    std_logic;
    spcptr0         : out    std_logic;
    spcptr1         : out    std_logic;
    spcptr2         : out    std_logic;
    spcptr3         : out    std_logic;
    spcptr4         : out    std_logic
  );
end entity;
