library ieee;
use ieee.std_logic_1164.all;

entity cadr_dram2 is
  port (
    dadr10c     : out std_logic;
    \-dadr0c\   : out std_logic;
    \-dadr1c\   : out std_logic;
    \-dadr2c\   : out std_logic;
    \-dadr3c\   : out std_logic;
    \-dadr4c\   : out std_logic;
    dpar        : out std_logic;
    \-dadr5c\   : out std_logic;
    \-dadr6c\   : out std_logic;
    \-dadr7c\   : out std_logic;
    \-dadr8c\   : out std_logic;
    \-dadr9c\   : out std_logic;
    \-dwec\     : out std_logic;
    aa17        : in  std_logic;
    \-dadr10c\  : out std_logic;
    dr          : out std_logic;
    aa16        : in  std_logic;
    r3          : in  std_logic;
    ir18b       : in  std_logic;
    hi11        : in  std_logic;
    dmask6      : in  std_logic;
    r6          : in  std_logic;
    ir15b       : in  std_logic;
    dmask3      : in  std_logic;
    dp          : out std_logic;
    aa15        : in  std_logic;
    dn          : out std_logic;
    aa14        : in  std_logic;
    r2          : in  std_logic;
    ir17b       : in  std_logic;
    dmask5      : in  std_logic;
    r5          : in  std_logic;
    ir14b       : in  std_logic;
    dmask2      : in  std_logic;
    dpc13       : out std_logic;
    aa13        : in  std_logic;
    dpc12       : out std_logic;
    aa12        : in  std_logic;
    r1          : in  std_logic;
    ir16b       : in  std_logic;
    dmask4      : in  std_logic;
    r4          : in  std_logic;
    ir13b       : in  std_logic;
    dmask1      : in  std_logic;
    ir12b       : in  std_logic;
    vmo19       : in  std_logic;
    ir9b        : in  std_logic;
    r0          : in  std_logic;
    dmask0      : in  std_logic;
    \-dmapbenb\ : in  std_logic;
    vmo18       : in  std_logic;
    ir8b        : in  std_logic;
    hi6         : in  std_logic;
    ir22b       : in  std_logic;
    ir21b       : in  std_logic;
    ir20b       : in  std_logic;
    ir19b       : in  std_logic;
    dispwr      : in  std_logic;
    wp2         : in  std_logic);
end;
