library ieee;
use ieee.std_logic_1164.all;

entity cadr_mctl is
  port (
    \-ir31\         : in     std_logic;
    clk4e           : in     std_logic;
    destmd          : in     std_logic;
    hi2             : in     std_logic;
    ir26            : in     std_logic;
    ir27            : in     std_logic;
    ir28            : in     std_logic;
    ir29            : in     std_logic;
    ir30            : in     std_logic;
    tse4a           : in     std_logic;
    wadr0           : in     std_logic;
    wadr1           : in     std_logic;
    wadr2           : in     std_logic;
    wadr3           : in     std_logic;
    wadr4           : in     std_logic;
    wp4b            : in     std_logic;
    \-madr0a\       : out    std_logic;
    \-madr0b\       : out    std_logic;
    \-madr1a\       : out    std_logic;
    \-madr1b\       : out    std_logic;
    \-madr2a\       : out    std_logic;
    \-madr2b\       : out    std_logic;
    \-madr3a\       : out    std_logic;
    \-madr3b\       : out    std_logic;
    \-madr4a\       : out    std_logic;
    \-madr4b\       : out    std_logic;
    \-mpass\        : out    std_logic;
    \-mpassl\       : out    std_logic;
    \-mpassm\       : out    std_logic;
    \-mwpa\         : out    std_logic;
    \-mwpb\         : out    std_logic;
    mmem0           : out    std_logic;
    mmem1           : out    std_logic;
    mmem10          : out    std_logic;
    mmem11          : out    std_logic;
    mmem12          : out    std_logic;
    mmem13          : out    std_logic;
    mmem14          : out    std_logic;
    mmem15          : out    std_logic;
    mmem16          : out    std_logic;
    mmem17          : out    std_logic;
    mmem18          : out    std_logic;
    mmem19          : out    std_logic;
    mmem2           : out    std_logic;
    mmem20          : out    std_logic;
    mmem21          : out    std_logic;
    mmem22          : out    std_logic;
    mmem23          : out    std_logic;
    mmem24          : out    std_logic;
    mmem25          : out    std_logic;
    mmem26          : out    std_logic;
    mmem27          : out    std_logic;
    mmem28          : out    std_logic;
    mmem29          : out    std_logic;
    mmem3           : out    std_logic;
    mmem30          : out    std_logic;
    mmem31          : out    std_logic;
    mmem4           : out    std_logic;
    mmem5           : out    std_logic;
    mmem6           : out    std_logic;
    mmem7           : out    std_logic;
    mmem8           : out    std_logic;
    mmem9           : out    std_logic;
    mmemparity      : out    std_logic;
    mpass           : out    std_logic;
    mpassl          : out    std_logic;
    srcm            : out    std_logic
  );
end entity cadr_mctl;
