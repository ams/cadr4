library ieee;
use ieee.std_logic_1164.all;

entity busint_lmadr is
  port (
    \-adr0\         : in     std_logic;
    \-adr10\        : in     std_logic;
    \-adr11\        : in     std_logic;
    \-adr12\        : in     std_logic;
    \-adr13\        : in     std_logic;
    \-adr14\        : in     std_logic;
    \-adr15\        : in     std_logic;
    \-adr16\        : in     std_logic;
    \-adr17\        : in     std_logic;
    \-adr18\        : in     std_logic;
    \-adr19\        : in     std_logic;
    \-adr1\         : in     std_logic;
    \-adr2\         : in     std_logic;
    \-adr3\         : in     std_logic;
    \-adr4\         : in     std_logic;
    \-adr5\         : in     std_logic;
    \-adr6\         : in     std_logic;
    \-adr7\         : in     std_logic;
    \-adr8\         : in     std_logic;
    \-adr9\         : in     std_logic;
    \-lmadr>ub\     : in     std_logic;
    \-lmadr>xbus\   : in     std_logic;
    uao1            : out    std_logic;
    uao10           : out    std_logic;
    uao11           : out    std_logic;
    uao12           : out    std_logic;
    uao13           : out    std_logic;
    uao14           : out    std_logic;
    uao15           : out    std_logic;
    uao16           : out    std_logic;
    uao17           : out    std_logic;
    uao2            : out    std_logic;
    uao3            : out    std_logic;
    uao4            : out    std_logic;
    uao5            : out    std_logic;
    uao6            : out    std_logic;
    uao7            : out    std_logic;
    uao8            : out    std_logic;
    uao9            : out    std_logic;
    xao0            : out    std_logic;
    xao1            : out    std_logic;
    xao10           : out    std_logic;
    xao11           : out    std_logic;
    xao12           : out    std_logic;
    xao13           : out    std_logic;
    xao14           : out    std_logic;
    xao15           : out    std_logic;
    xao16           : out    std_logic;
    xao17           : out    std_logic;
    xao18           : out    std_logic;
    xao19           : out    std_logic;
    xao2            : out    std_logic;
    xao3            : out    std_logic;
    xao4            : out    std_logic;
    xao5            : out    std_logic;
    xao6            : out    std_logic;
    xao7            : out    std_logic;
    xao8            : out    std_logic;
    xao9            : out    std_logic
  );
end entity;
