library ieee;
use ieee.std_logic_1164.all;

entity busint_xd is
  port (
    \-xdrive\       : in     std_logic;
    \hi 15-30\      : in     std_logic;
    \xbus par out\  : in     std_logic;
    bus0            : in     std_logic;
    bus1            : in     std_logic;
    bus10           : in     std_logic;
    bus11           : in     std_logic;
    bus12           : in     std_logic;
    bus13           : in     std_logic;
    bus14           : in     std_logic;
    bus15           : in     std_logic;
    bus16           : in     std_logic;
    bus17           : in     std_logic;
    bus18           : in     std_logic;
    bus19           : in     std_logic;
    bus2            : in     std_logic;
    bus20           : in     std_logic;
    bus21           : in     std_logic;
    bus22           : in     std_logic;
    bus23           : in     std_logic;
    bus24           : in     std_logic;
    bus25           : in     std_logic;
    bus26           : in     std_logic;
    bus27           : in     std_logic;
    bus28           : in     std_logic;
    bus29           : in     std_logic;
    bus3            : in     std_logic;
    bus30           : in     std_logic;
    bus31           : in     std_logic;
    bus4            : in     std_logic;
    bus5            : in     std_logic;
    bus6            : in     std_logic;
    bus7            : in     std_logic;
    bus8            : in     std_logic;
    bus9            : in     std_logic;
    \-xbus ignpar\  : inout  std_logic;
    \-xbus par\     : inout  std_logic;
    \-xbus wr\      : inout  std_logic;
    \-xbus0\        : inout  std_logic;
    \-xbus10\       : inout  std_logic;
    \-xbus11\       : inout  std_logic;
    \-xbus12\       : inout  std_logic;
    \-xbus13\       : inout  std_logic;
    \-xbus14\       : inout  std_logic;
    \-xbus15\       : inout  std_logic;
    \-xbus16\       : inout  std_logic;
    \-xbus17\       : inout  std_logic;
    \-xbus18\       : inout  std_logic;
    \-xbus19\       : inout  std_logic;
    \-xbus1\        : inout  std_logic;
    \-xbus20\       : inout  std_logic;
    \-xbus21\       : inout  std_logic;
    \-xbus22\       : inout  std_logic;
    \-xbus23\       : inout  std_logic;
    \-xbus24\       : inout  std_logic;
    \-xbus25\       : inout  std_logic;
    \-xbus26\       : inout  std_logic;
    \-xbus27\       : inout  std_logic;
    \-xbus28\       : inout  std_logic;
    \-xbus29\       : inout  std_logic;
    \-xbus2\        : inout  std_logic;
    \-xbus30\       : inout  std_logic;
    \-xbus31\       : inout  std_logic;
    \-xbus3\        : inout  std_logic;
    \-xbus4\        : inout  std_logic;
    \-xbus5\        : inout  std_logic;
    \-xbus6\        : inout  std_logic;
    \-xbus7\        : inout  std_logic;
    \-xbus8\        : inout  std_logic;
    \-xbus9\        : inout  std_logic;
    \xbus ignpar in\ : out    std_logic;
    \xbus par in\   : out    std_logic;
    xdi0            : out    std_logic;
    xdi1            : out    std_logic;
    xdi10           : out    std_logic;
    xdi11           : out    std_logic;
    xdi12           : out    std_logic;
    xdi13           : out    std_logic;
    xdi14           : out    std_logic;
    xdi15           : out    std_logic;
    xdi16           : out    std_logic;
    xdi17           : out    std_logic;
    xdi18           : out    std_logic;
    xdi19           : out    std_logic;
    xdi2            : out    std_logic;
    xdi20           : out    std_logic;
    xdi21           : out    std_logic;
    xdi22           : out    std_logic;
    xdi23           : out    std_logic;
    xdi24           : out    std_logic;
    xdi25           : out    std_logic;
    xdi26           : out    std_logic;
    xdi27           : out    std_logic;
    xdi28           : out    std_logic;
    xdi29           : out    std_logic;
    xdi3            : out    std_logic;
    xdi30           : out    std_logic;
    xdi31           : out    std_logic;
    xdi4            : out    std_logic;
    xdi5            : out    std_logic;
    xdi6            : out    std_logic;
    xdi7            : out    std_logic;
    xdi8            : out    std_logic;
    xdi9            : out    std_logic
  );
end entity;
