library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_7464 is
  port (
    d4    : in  std_logic;
    b2    : in  std_logic;
    a2    : in  std_logic;
    c3    : in  std_logic;
    b3    : in  std_logic;
    a3    : in  std_logic;
    \out\ : out std_logic;
    a1    : in  std_logic;
    b1    : in  std_logic;
    c4    : in  std_logic;
    b4    : in  std_logic;
    a4    : in  std_logic
    );
end ic_7464;

architecture ttl of ic_7464 is
begin

end ttl;
