library ieee;
use ieee.std_logic_1164.all;

entity icmem_olord2 is
  port (
    \-busint.lm.reset\ : in     std_logic;
    \-halt\         : in     std_logic;
    \-ldmode\       : in     std_logic;
    \-upperhighok\  : in     std_logic;
    \prog.bus.reset\ : in     std_logic;
    \stat.ovf\      : in     std_logic;
    aparok          : in     std_logic;
    clk5            : in     std_logic;
    dparok          : in     std_logic;
    errstop         : in     std_logic;
    iparok          : in     std_logic;
    mclk5           : in     std_logic;
    memparok        : in     std_logic;
    mmemparok       : in     std_logic;
    pdlparok        : in     std_logic;
    spcparok        : in     std_logic;
    spy6            : in     std_logic;
    spy7            : in     std_logic;
    srun            : in     std_logic;
    v0parok         : in     std_logic;
    vmoparok        : in     std_logic;
    \-ape\          : out    std_logic;
    \-boot1\        : out    std_logic;
    \-boot2\        : out    std_logic;
    \-boot\         : out    std_logic;
    \-bus.power.reset\ : out    std_logic;
    \-bus.reset\    : out    std_logic;
    \-clk5\         : out    std_logic;
    \-clock reset a\ : out    std_logic;
    \-clock reset b\ : out    std_logic;
    \-dpe\          : out    std_logic;
    \-errhalt\      : out    std_logic;
    \-halted\       : out    std_logic;
    \-higherr\      : out    std_logic;
    \-ipe\          : out    std_logic;
    \-lowerhighok\  : out    std_logic;
    \-mclk5\        : out    std_logic;
    \-mempe\        : out    std_logic;
    \-mpe\          : out    std_logic;
    \-pdlpe\        : out    std_logic;
    \-power reset\  : out    std_logic;
    \-prog.reset\   : out    std_logic;
    \-reset\        : out    std_logic;
    \-spe\          : out    std_logic;
    \-v0pe\         : out    std_logic;
    \-v1pe\         : out    std_logic;
    \boot.trap\     : out    std_logic;
    \power reset a\ : out    std_logic;
    \prog.boot\     : out    std_logic;
    clk5a           : out    std_logic;
    err             : out    std_logic;
    hi1             : out    std_logic;
    hi2             : out    std_logic;
    highok          : out    std_logic;
    ldmode          : out    std_logic;
    mclk5a          : out    std_logic;
    reset           : out    std_logic;
    statstop        : out    std_logic
  );
end entity;
