library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_vma is
  port (
    \-vmadrive\ : out std_logic;
    \-vma31\    : out std_logic;
    mf24        : out std_logic;
    \-vma30\    : out std_logic;
    mf25        : out std_logic;
    \-vma29\    : out std_logic;
    mf26        : out std_logic;
    \-vma28\    : out std_logic;
    mf27        : out std_logic;
    \-vma27\    : out std_logic;
    mf28        : out std_logic;
    \-vma26\    : out std_logic;
    mf29        : out std_logic;
    \-vma25\    : out std_logic;
    mf30        : out std_logic;
    \-vma24\    : out std_logic;
    mf31        : out std_logic;
    \-vma7\     : out std_logic;
    mf0         : out std_logic;
    \-vma6\     : out std_logic;
    mf1         : out std_logic;
    \-vma5\     : out std_logic;
    mf2         : out std_logic;
    \-vma4\     : out std_logic;
    mf3         : out std_logic;
    \-vma3\     : out std_logic;
    mf4         : out std_logic;
    \-vma2\     : out std_logic;
    mf5         : out std_logic;
    \-vma1\     : out std_logic;
    mf6         : out std_logic;
    \-vma0\     : out std_logic;
    mf7         : out std_logic;
    \-vma23\    : out std_logic;
    mf16        : out std_logic;
    \-vma22\    : out std_logic;
    mf17        : out std_logic;
    \-vma21\    : out std_logic;
    mf18        : out std_logic;
    \-vma20\    : out std_logic;
    mf19        : out std_logic;
    \-vma19\    : out std_logic;
    mf20        : out std_logic;
    \-vma18\    : out std_logic;
    mf21        : out std_logic;
    \-vma17\    : out std_logic;
    mf22        : out std_logic;
    \-vma16\    : out std_logic;
    mf23        : out std_logic;
    \-vma15\    : out std_logic;
    mf8         : out std_logic;
    \-vma14\    : out std_logic;
    mf9         : out std_logic;
    \-vma13\    : out std_logic;
    mf10        : out std_logic;
    \-vma12\    : out std_logic;
    mf11        : out std_logic;
    \-vma11\    : out std_logic;
    mf12        : out std_logic;
    \-vma10\    : out std_logic;
    mf13        : out std_logic;
    \-vma9\     : out std_logic;
    mf14        : out std_logic;
    \-vma8\     : out std_logic;
    mf15        : out std_logic;
    tse2        : in  std_logic;
    srcvma      : out std_logic;
    \-vmaenb\   : in  std_logic;
    \-vmas24\   : in  std_logic;
    \-vmas25\   : in  std_logic;
    \-vmas26\   : in  std_logic;
    clk1a       : in  std_logic;
    \-vmas27\   : in  std_logic;
    \-vmas28\   : in  std_logic;
    \-vmas29\   : in  std_logic;
    \-vmas30\   : in  std_logic;
    \-vmas31\   : in  std_logic;
    \-vmas0\    : in  std_logic;
    \-vmas1\    : in  std_logic;
    \-vmas2\    : in  std_logic;
    clk2a       : in  std_logic;
    \-vmas3\    : in  std_logic;
    \-vmas4\    : in  std_logic;
    \-vmas5\    : in  std_logic;
    \-vmas12\   : in  std_logic;
    \-vmas13\   : in  std_logic;
    \-vmas14\   : in  std_logic;
    \-vmas15\   : in  std_logic;
    \-vmas16\   : in  std_logic;
    \-vmas17\   : in  std_logic;
    \-vmas18\   : in  std_logic;
    \-vmas19\   : in  std_logic;
    \-vmas20\   : in  std_logic;
    \-vmas21\   : in  std_logic;
    \-vmas22\   : in  std_logic;
    \-vmas23\   : in  std_logic;
    \-vmas6\    : in  std_logic;
    \-vmas7\    : in  std_logic;
    \-vmas8\    : in  std_logic;
    clk2c       : in  std_logic;
    \-vmas9\    : in  std_logic;
    \-vmas10\   : in  std_logic;
    \-vmas11\   : in  std_logic;
    \-srcvma\   : in  std_logic);
end;

architecture ttl of cadr_vma is
  signal nc115 : std_logic;
  signal nc116 : std_logic;
  signal nc117 : std_logic;
  signal nc118 : std_logic;
  signal nc119 : std_logic;
  signal nc120 : std_logic;
  signal nc121 : std_logic;
  signal nc122 : std_logic;
begin
  vma_1a06 : sn74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma31\, bout3 => mf24, ain1 => \-vma30\, bout2 => mf25, ain2 => \-vma29\, bout1 => mf26, ain3 => \-vma28\, bout0 => mf27, bin0 => \-vma27\, aout3 => mf28, bin1 => \-vma26\, aout2 => mf29, bin2 => \-vma25\, aout1 => mf30, bin3 => \-vma24\, aout0 => mf31, benb_n => \-vmadrive\);
  vma_1a10 : sn74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma7\, bout3 => mf0, ain1 => \-vma6\, bout2 => mf1, ain2 => \-vma5\, bout1 => mf2, ain3 => \-vma4\, bout0 => mf3, bin0 => \-vma3\, aout3 => mf4, bin1 => \-vma2\, aout2 => mf5, bin2 => \-vma1\, aout1 => mf6, bin3 => \-vma0\, aout0 => mf7, benb_n => \-vmadrive\);
  vma_1a12 : sn74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma23\, bout3 => mf16, ain1 => \-vma22\, bout2 => mf17, ain2 => \-vma21\, bout1 => mf18, ain3 => \-vma20\, bout0 => mf19, bin0 => \-vma19\, aout3 => mf20, bin1 => \-vma18\, aout2 => mf21, bin2 => \-vma17\, aout1 => mf22, bin3 => \-vma16\, aout0 => mf23, benb_n => \-vmadrive\);
  vma_1a14 : sn74s240 port map(aenb_n => \-vmadrive\, ain0 => \-vma15\, bout3 => mf8, ain1 => \-vma14\, bout2 => mf9, ain2 => \-vma13\, bout1 => mf10, ain3 => \-vma12\, bout0 => mf11, bin0 => \-vma11\, aout3 => mf12, bin1 => \-vma10\, aout2 => mf13, bin2 => \-vma9\, aout1 => mf14, bin3 => \-vma8\, aout0 => mf15, benb_n => \-vmadrive\);
  vma_1a18 : sn74s00 port map(g4q_n   => \-vmadrive\, g4a => tse2, g4b => srcvma, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3b => '0', g3a => '0');
  vma_1b22 : am25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma24\, i0 => \-vmas24\, i1 => \-vmas25\, d1 => \-vma25\, i2 => \-vmas26\, d2 => \-vma26\, clk => clk1a, d3 => \-vma27\, i3 => \-vmas27\, d4 => \-vma28\, i4 => \-vmas28\, i5 => \-vmas29\, d5 => \-vma29\);
  vma_1b23 : am25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma30\, i0 => \-vmas30\, i1 => \-vmas31\, d1 => \-vma31\, i2 => nc115, d2 => nc116, clk => clk1a, d3 => nc117, i3 => nc118, d4 => nc119, i4 => nc120, i5 => nc121, d5 => nc122);
  vma_1c22 : am25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma0\, i0 => \-vmas0\, i1 => \-vmas1\, d1 => \-vma1\, i2 => \-vmas2\, d2 => \-vma2\, clk => clk2a, d3 => \-vma3\, i3 => \-vmas3\, d4 => \-vma4\, i4 => \-vmas4\, i5 => \-vmas5\, d5 => \-vma5\);
  vma_1c24 : am25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma12\, i0 => \-vmas12\, i1 => \-vmas13\, d1 => \-vma13\, i2 => \-vmas14\, d2 => \-vma14\, clk => clk2a, d3 => \-vma15\, i3 => \-vmas15\, d4 => \-vma16\, i4 => \-vmas16\, i5 => \-vmas17\, d5 => \-vma17\);
  vma_1c25 : am25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma18\, i0 => \-vmas18\, i1 => \-vmas19\, d1 => \-vma19\, i2 => \-vmas20\, d2 => \-vma20\, clk => clk2a, d3 => \-vma21\, i3 => \-vmas21\, d4 => \-vma22\, i4 => \-vmas22\, i5 => \-vmas23\, d5 => \-vma23\);
  vma_1d25 : am25s07 port map(enb_n   => \-vmaenb\, d0 => \-vma6\, i0 => \-vmas6\, i1 => \-vmas7\, d1 => \-vma7\, i2 => \-vmas8\, d2 => \-vma8\, clk => clk2c, d3 => \-vma9\, i3 => \-vmas9\, d4 => \-vma10\, i4 => \-vmas10\, i5 => \-vmas11\, d5 => \-vma11\);
  vma_2a05 : sn74s04 port map(g3a     => \-srcvma\, g3q_n => srcvma, g1a => '0', g2a => '0', g4a => '0', g5a => '0', g6a => '0');
end architecture;
