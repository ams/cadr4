library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_7451 is
  port (
    g1a : in  std_logic;
    g2a : in  std_logic;
    g2b : in  std_logic;
    g2c : in  std_logic;
    g2d : in  std_logic;
    g2y : out std_logic;
    g1y : out std_logic;
    g1c : in  std_logic;
    g1d : in  std_logic;
    g1b : in  std_logic
    );
end ic_7451;

architecture ttl of ic_7451 is
begin

end ttl;
