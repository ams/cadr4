library ieee;
use ieee.std_logic_1164.all;

entity cadr_source is
  port (
    \-idebug\       : in     std_logic;
    \-ir31\         : in     std_logic;
    \-iwrited\      : in     std_logic;
    hi5             : in     std_logic;
    ir10            : in     std_logic;
    ir11            : in     std_logic;
    ir19            : in     std_logic;
    ir20            : in     std_logic;
    ir21            : in     std_logic;
    ir22            : in     std_logic;
    ir23            : in     std_logic;
    ir25            : in     std_logic;
    ir26            : in     std_logic;
    ir27            : in     std_logic;
    ir28            : in     std_logic;
    ir29            : in     std_logic;
    ir3             : in     std_logic;
    ir4             : in     std_logic;
    ir43            : in     std_logic;
    ir44            : in     std_logic;
    ir8             : in     std_logic;
    nop             : in     std_logic;
    \-destimod0\    : out    std_logic;
    \-destimod1\    : out    std_logic;
    \-destintctl\   : out    std_logic;
    \-destlc\       : out    std_logic;
    \-destmdr\      : out    std_logic;
    \-destmem\      : out    std_logic;
    \-destpdl(p)\   : out    std_logic;
    \-destpdl(x)\   : out    std_logic;
    \-destpdlp\     : out    std_logic;
    \-destpdltop\   : out    std_logic;
    \-destpdlx\     : out    std_logic;
    \-destspc\      : out    std_logic;
    \-destvma\      : out    std_logic;
    \-div\          : out    std_logic;
    \-funct0\       : out    std_logic;
    \-funct1\       : out    std_logic;
    \-funct2\       : out    std_logic;
    \-funct3\       : out    std_logic;
    \-ir22\         : out    std_logic;
    \-ir25\         : out    std_logic;
    \-iralu\        : out    std_logic;
    \-irbyte\       : out    std_logic;
    \-irdisp\       : out    std_logic;
    \-irjump\       : out    std_logic;
    \-mul\          : out    std_logic;
    \-specalu\      : out    std_logic;
    \-srcdc\        : out    std_logic;
    \-srclc\        : out    std_logic;
    \-srcmap\       : out    std_logic;
    \-srcmd\        : out    std_logic;
    \-srcopc\       : out    std_logic;
    \-srcpdlidx\    : out    std_logic;
    \-srcpdlpop\    : out    std_logic;
    \-srcpdlptr\    : out    std_logic;
    \-srcpdltop\    : out    std_logic;
    \-srcq\         : out    std_logic;
    \-srcspc\       : out    std_logic;
    \-srcspcpop\    : out    std_logic;
    \-srcvma\       : out    std_logic;
    dest            : out    std_logic;
    destm           : out    std_logic;
    imod            : out    std_logic;
    iralu           : out    std_logic;
    irdisp          : out    std_logic;
    irjump          : out    std_logic
  );
end entity cadr_source;
