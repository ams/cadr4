library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_vmem1 is
  port (
    \-vma17\   : in  std_logic;
    \-vma18\   : in  std_logic;
    \-vma19\   : in  std_logic;
    \-vma20\   : in  std_logic;
    \-vma21\   : in  std_logic;
    \-vma22\   : in  std_logic;
    \-vma23\   : in  std_logic;
    vm1mpar    : out std_logic;
    \-vma12\   : in  std_logic;
    \-vma13\   : in  std_logic;
    \-vma14\   : in  std_logic;
    \-vma15\   : in  std_logic;
    \-vma16\   : in  std_logic;
    \-vma5\    : in  std_logic;
    \-vma6\    : in  std_logic;
    \-vma7\    : in  std_logic;
    \-vma8\    : in  std_logic;
    \-vma9\    : in  std_logic;
    \-vma10\   : in  std_logic;
    \-vma11\   : in  std_logic;
    \-vm1lpar\ : out std_logic;
    \-vma0\    : in  std_logic;
    \-vma1\    : in  std_logic;
    \-vma2\    : in  std_logic;
    \-vma3\    : in  std_logic;
    \-vma4\    : in  std_logic;
    gnd        : in  std_logic;
    vmap4a     : out std_logic;
    vmap3a     : out std_logic;
    vmap2a     : out std_logic;
    vmap1a     : out std_logic;
    vmap0a     : out std_logic;
    \-vmo10\   : out std_logic;
    \-mapi12a\ : out std_logic;
    \-mapi11a\ : out std_logic;
    \-mapi10a\ : out std_logic;
    \-mapi9a\  : out std_logic;
    \-mapi8a\  : out std_logic;
    \-vm1wpa\  : in  std_logic;
    \-vmo4\    : out std_logic;
    \-vmo2\    : out std_logic;
    mapi10     : in  std_logic;
    mapi9      : in  std_logic;
    mapi8      : in  std_logic;
    \-vmap4\   : in  std_logic;
    \-vmap3\   : in  std_logic;
    \-vmap2\   : in  std_logic;
    \-vmap1\   : in  std_logic;
    \-vmap0\   : in  std_logic;
    \-vmo0\    : out std_logic;
    vm1pari    : out std_logic;
    mapi12     : in  std_logic;
    mapi11     : in  std_logic;
    \-mapi8b\  : out std_logic;
    \-mapi9b\  : out std_logic;
    \-mapi10b\ : out std_logic;
    \-mapi11b\ : out std_logic;
    \-mapi12b\ : out std_logic;
    \-vmo11\   : out std_logic;
    \-vmo5\    : out std_logic;
    \-vmo9\    : out std_logic;
    \-vmo3\    : out std_logic;
    \-vmo8\    : out std_logic;
    \-vmo7\    : out std_logic;
    \-vmo1\    : out std_logic;
    \-vmo6\    : out std_logic);
end;

architecture ttl of cadr_vmem1 is
  signal nc109 : std_logic;
  signal nc110 : std_logic;
  signal nc111 : std_logic;
  signal nc112 : std_logic;
begin
  vmem1_1c03 : am93s48 port map(i6      => \-vma17\, i5 => \-vma18\, i4 => \-vma19\, i3 => \-vma20\, i2 => \-vma21\, i1 => \-vma22\, i0 => \-vma23\, po => vm1mpar, pe => nc109, i11 => \-vma12\, i10 => \-vma13\, i9 => \-vma14\, i8 => \-vma15\, i7 => \-vma16\);
  vmem1_1c04 : am93s48 port map(i6      => \-vma5\, i5 => \-vma6\, i4 => \-vma7\, i3 => \-vma8\, i2 => \-vma9\, i1 => \-vma10\, i0 => \-vma11\, po => nc110, pe => \-vm1lpar\, i11 => \-vma0\, i10 => \-vma1\, i9 => \-vma2\, i8 => \-vma3\, i7 => \-vma4\);
  vmem1_1d01 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo10\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma10\);
  vmem1_1d02 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo4\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma4\);
  vmem1_1d06 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo2\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma2\);
  vmem1_1d08 : sn74s240 port map(aenb_n => gnd, ain0 => mapi10, bout3 => vmap0a, ain1 => mapi9, bout2 => vmap1a, ain2 => mapi8, bout1 => vmap2a, ain3 => \-vmap4\, bout0 => vmap3a, bin0 => \-vmap3\, aout3 => vmap4a, bin1 => \-vmap2\, aout2 => \-mapi8a\, bin2 => \-vmap1\, aout1 => \-mapi9a\, bin3 => \-vmap0\, aout0 => \-mapi10a\, benb_n => gnd);
  vmem1_1d11 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo0\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma0\);
  vmem1_1d12 : sn74s86 port map(g1a     => vm1mpar, g1b => \-vm1lpar\, g1y => vm1pari, g2a => '0', g2b => '0', g3a => '0', g3b => '0', g4a => '0', g4b => '0');
  vmem1_1d13 : sn74s240 port map(aenb_n => gnd, ain0 => mapi12, bout3 => \-mapi11a\, ain1 => mapi11, bout2 => \-mapi12a\, ain2 => mapi10, bout1 => nc111, ain3 => mapi9, bout0 => \-mapi8b\, bin0 => mapi8, aout3 => \-mapi9b\, bin1 => nc112, aout2 => \-mapi10b\, bin2 => mapi12, aout1 => \-mapi11b\, bin3 => mapi11, aout0 => \-mapi12b\, benb_n => gnd);
  vmem1_1e04 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo11\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma11\);
  vmem1_1e05 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo5\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma5\);
  vmem1_1e08 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo9\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma9\);
  vmem1_1e09 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo3\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma3\);
  vmem1_1e10 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo8\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma8\);
  vmem1_1e13 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo7\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma7\);
  vmem1_1e14 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo1\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma1\);
  vmem1_1e15 : am93425a port map(ce_n   => gnd, a0 => vmap4a, a1 => vmap3a, a2 => vmap2a, a3 => vmap1a, a4 => vmap0a, do => \-vmo6\, a5 => \-mapi12a\, a6 => \-mapi11a\, a7 => \-mapi10a\, a8 => \-mapi9a\, a9 => \-mapi8a\, we_n => \-vm1wpa\, di => \-vma6\);
end architecture;
