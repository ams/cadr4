library ieee;
use ieee.std_logic_1164.all;

entity icmem_stat is
  port (
    \-ldstat\       : in     std_logic;
    \-spy.sth\      : in     std_logic;
    \-spy.stl\      : in     std_logic;
    \-statbit\      : in     std_logic;
    clk5a           : in     std_logic;
    hi1             : in     std_logic;
    iwr0            : in     std_logic;
    iwr1            : in     std_logic;
    iwr10           : in     std_logic;
    iwr11           : in     std_logic;
    iwr12           : in     std_logic;
    iwr13           : in     std_logic;
    iwr14           : in     std_logic;
    iwr15           : in     std_logic;
    iwr16           : in     std_logic;
    iwr17           : in     std_logic;
    iwr18           : in     std_logic;
    iwr19           : in     std_logic;
    iwr2            : in     std_logic;
    iwr20           : in     std_logic;
    iwr21           : in     std_logic;
    iwr22           : in     std_logic;
    iwr23           : in     std_logic;
    iwr24           : in     std_logic;
    iwr25           : in     std_logic;
    iwr26           : in     std_logic;
    iwr27           : in     std_logic;
    iwr28           : in     std_logic;
    iwr29           : in     std_logic;
    iwr3            : in     std_logic;
    iwr30           : in     std_logic;
    iwr31           : in     std_logic;
    iwr4            : in     std_logic;
    iwr5            : in     std_logic;
    iwr6            : in     std_logic;
    iwr7            : in     std_logic;
    iwr8            : in     std_logic;
    iwr9            : in     std_logic;
    \-stc12\        : out    std_logic;
    \-stc16\        : out    std_logic;
    \-stc20\        : out    std_logic;
    \-stc24\        : out    std_logic;
    \-stc28\        : out    std_logic;
    \-stc32\        : out    std_logic;
    \-stc4\         : out    std_logic;
    \-stc8\         : out    std_logic;
    spy0            : out    std_logic;
    spy1            : out    std_logic;
    spy10           : out    std_logic;
    spy11           : out    std_logic;
    spy12           : out    std_logic;
    spy13           : out    std_logic;
    spy14           : out    std_logic;
    spy15           : out    std_logic;
    spy2            : out    std_logic;
    spy3            : out    std_logic;
    spy4            : out    std_logic;
    spy5            : out    std_logic;
    spy6            : out    std_logic;
    spy7            : out    std_logic;
    spy8            : out    std_logic;
    spy9            : out    std_logic;
    st0             : out    std_logic;
    st1             : out    std_logic;
    st10            : out    std_logic;
    st11            : out    std_logic;
    st12            : out    std_logic;
    st13            : out    std_logic;
    st14            : out    std_logic;
    st15            : out    std_logic;
    st16            : out    std_logic;
    st17            : out    std_logic;
    st18            : out    std_logic;
    st19            : out    std_logic;
    st2             : out    std_logic;
    st20            : out    std_logic;
    st21            : out    std_logic;
    st22            : out    std_logic;
    st23            : out    std_logic;
    st24            : out    std_logic;
    st25            : out    std_logic;
    st26            : out    std_logic;
    st27            : out    std_logic;
    st28            : out    std_logic;
    st29            : out    std_logic;
    st3             : out    std_logic;
    st30            : out    std_logic;
    st31            : out    std_logic;
    st4             : out    std_logic;
    st5             : out    std_logic;
    st6             : out    std_logic;
    st7             : out    std_logic;
    st8             : out    std_logic;
    st9             : out    std_logic
  );
end entity;
