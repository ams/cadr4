library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr4;
use cadr4.utilities.all;

entity cadr4_clockd is
  port (
    \-clk1\        : out std_logic;
    hi12           : in  std_logic;
    clk1a          : out std_logic;
    reset          : in  std_logic;
    \-reset\       : out std_logic;
    mclk1a         : out std_logic;
    \-mclk1\       : out std_logic;
    mclk1          : in  std_logic;
    clk1           : in  std_logic;
    \-wp1\         : in  std_logic;
    wp1b           : out std_logic;
    wp1a           : out std_logic;
    tse1b          : out std_logic;
    \-tse1\        : in  std_logic;
    tse1a          : out std_logic;
    hi1            : in  std_logic;
    hi2            : in  std_logic;
    hi3            : in  std_logic;
    hi4            : in  std_logic;
    hi5            : in  std_logic;
    hi6            : in  std_logic;
    hi7            : in  std_logic;
    \-upperhighok\ : out std_logic;
    hi8            : in  std_logic;
    hi9            : in  std_logic;
    hi10           : in  std_logic;
    hi11           : in  std_logic;
    lcry3          : in  std_logic;
    \-lcry3\       : out std_logic;
    nc429          : in  std_logic;
    nc430          : out std_logic;
    clk2           : in  std_logic;
    \-clk2c\       : out std_logic;
    \-clk2a\       : out std_logic;
    wp2            : out std_logic;
    \-wp2\         : in  std_logic;
    tse2           : out std_logic;
    \-tse2\        : in  std_logic;
    clk2a          : out std_logic;
    clk2b          : out std_logic;
    clk2c          : out std_logic;
    \-clk3a\       : out std_logic;
    clk3a          : out std_logic;
    clk3b          : out std_logic;
    clk3c          : out std_logic;
    nc427          : in  std_logic;
    nc428          : out std_logic;
    clk3           : in  std_logic;
    \-clk3g\       : out std_logic;
    \-clk3d\       : out std_logic;
    wp3a           : out std_logic;
    \-wp3\         : in  std_logic;
    tse3a          : out std_logic;
    \-tse3\        : in  std_logic;
    clk3d          : out std_logic;
    clk3e          : out std_logic;
    clk3f          : out std_logic;
    \-clk4a\       : out std_logic;
    clk4a          : out std_logic;
    clk4b          : out std_logic;
    clk4c          : out std_logic;
    clk4           : in  std_logic;
    \-clk4e\       : out std_logic;
    \-clk4d\       : out std_logic;
    wp4c           : out std_logic;
    \-wp4\         : in  std_logic;
    wp4b           : out std_logic;
    wp4a           : out std_logic;
    clk4d          : out std_logic;
    clk4e          : out std_logic;
    clk4f          : out std_logic;
    nc423          : in  std_logic;
    nc424          : out std_logic;
    nc425          : in  std_logic;
    nc426          : out std_logic;
    \-tse4\        : in  std_logic;
    tse4b          : out std_logic;
    tse4a          : out std_logic;
    srcpdlptr      : out std_logic;
    \-srcpdlptr\   : in  std_logic;
    srcpdlidx      : out std_logic;
    \-srcpdlidx\   : in  std_logic);
end;

architecture ttl of cadr4_clockd is
begin
  clockd_1b18 : sn74s37 port map(g1a => \-clk1\, g1b => hi12, g1y => clk1a, g2a => reset, g2b => hi12, g2y => \-reset\, g3y => mclk1a, g3a => hi12, g3b => \-mclk1\, g4a => '0', g4b => '0');
  clockd_1b19 : sn74s04 port map(g1a => mclk1, g1q_n => \-mclk1\, g2a => clk1, g2q_n => \-clk1\, g3a => \-wp1\, g3q_n => wp1b, g4q_n => wp1a, g4a => \-wp1\, g5q_n => tse1b, g5a => \-tse1\, g6q_n => tse1a, g6a => \-tse1\);
  clockd_1f05 : sn74s133 port map(g  => hi1, f => hi2, e => hi3, d => hi4, c => hi5, b => hi6, a => hi7, q_n => \-upperhighok\, h => hi8, i => hi9, j => hi10, k => hi11, l => hi12, m => hi11);
  clockd_2c02 : sn74s04 port map(g1a => lcry3, g1q_n => \-lcry3\, g2a => nc429, g2q_n => nc430, g3a => clk2, g3q_n => \-clk2c\, g4q_n => \-clk2a\, g4a => clk2, g5q_n => wp2, g5a => \-wp2\, g6q_n => tse2, g6a => \-tse2\);
  clockd_2c03 : sn74s37 port map(g1a => \-clk2a\, g1b => hi7, g1y => clk2a, g2a => \-clk2a\, g2b => hi7, g2y => clk2b, g3y => clk2c, g3a => hi7, g3b => \-clk2c\, g4a => '0', g4b => '0');
  clockd_3c11 : sn74s37 port map(g1a => \-clk3a\, g1b => hi5, g1y => clk3a, g2a => \-clk3a\, g2b => hi5, g2y => clk3b, g3y => clk3c, g3a => hi5, g3b => \-clk3a\, g4a => '0', g4b => '0');
  clockd_3c12 : sn74s04 port map(g1a => nc427, g1q_n => nc428, g2a => clk3, g2q_n => \-clk3g\, g3a => clk3, g3q_n => \-clk3d\, g4q_n => \-clk3a\, g4a => clk3, g5q_n => wp3a, g5a => \-wp3\, g6q_n => tse3a, g6a => \-tse3\);
  clockd_3c13 : sn74s37 port map(g1a => \-clk3d\, g1b => hi5, g1y => clk3d, g2a => \-clk3d\, g2b => hi5, g2y => clk3e, g3y => clk3f, g3a => hi5, g3b => \-clk3d\, g4a => '0', g4b => '0');
  clockd_4c02 : sn74s37 port map(g1a => \-clk4a\, g1b => hi5, g1y => clk4a, g2a => \-clk4a\, g2b => hi5, g2y => clk4b, g3y => clk4c, g3a => hi5, g3b => \-clk4a\, g4a => '0', g4b => '0');
  clockd_4c06 : sn74s04 port map(g1a => clk4, g1q_n => \-clk4e\, g2a => clk4, g2q_n => \-clk4d\, g3a => clk4, g3q_n => \-clk4a\, g4q_n => wp4c, g4a => \-wp4\, g5q_n => wp4b, g5a => \-wp4\, g6q_n => wp4a, g6a => \-wp4\);
  clockd_4c07 : sn74s37 port map(g1a => \-clk4d\, g1b => hi2, g1y => clk4d, g2a => \-clk4d\, g2b => hi2, g2y => clk4e, g3y => clk4f, g3a => hi2, g3b => \-clk4d\, g4a => '0', g4b => '0');
  clockd_4d03 : sn74s04 port map(g1a => nc423, g1q_n => nc424, g2a => nc425, g2q_n => nc426, g3a => \-tse4\, g3q_n => tse4b, g4q_n => tse4a, g4a => \-tse4\, g5q_n => srcpdlptr, g5a => \-srcpdlptr\, g6q_n => srcpdlidx, g6a => \-srcpdlidx\);
end architecture;
