library ieee;
use ieee.std_logic_1164.all;

entity cadr_l is
  port (
    l7         : out std_logic;
    ob7        : in  std_logic;
    ob6        : in  std_logic;
    l6         : out std_logic;
    l5         : out std_logic;
    ob5        : in  std_logic;
    ob4        : in  std_logic;
    l4         : out std_logic;
    clk3f      : in  std_logic;
    l3         : out std_logic;
    ob3        : in  std_logic;
    ob2        : in  std_logic;
    l2         : out std_logic;
    l1         : out std_logic;
    ob1        : in  std_logic;
    ob0        : in  std_logic;
    l0         : out std_logic;
    l15        : out std_logic;
    ob15       : in  std_logic;
    ob14       : in  std_logic;
    l14        : out std_logic;
    l13        : out std_logic;
    ob13       : in  std_logic;
    ob12       : in  std_logic;
    l12        : out std_logic;
    l11        : out std_logic;
    ob11       : in  std_logic;
    ob10       : in  std_logic;
    l10        : out std_logic;
    l9         : out std_logic;
    ob9        : in  std_logic;
    ob8        : in  std_logic;
    l8         : out std_logic;
    l23        : out std_logic;
    ob23       : in  std_logic;
    ob22       : in  std_logic;
    l22        : out std_logic;
    l21        : out std_logic;
    ob21       : in  std_logic;
    ob20       : in  std_logic;
    l20        : out std_logic;
    l19        : out std_logic;
    ob19       : in  std_logic;
    ob18       : in  std_logic;
    l18        : out std_logic;
    l17        : out std_logic;
    ob17       : in  std_logic;
    ob16       : in  std_logic;
    l16        : out std_logic;
    l31        : out std_logic;
    ob31       : in  std_logic;
    ob30       : in  std_logic;
    l30        : out std_logic;
    l29        : out std_logic;
    ob29       : in  std_logic;
    ob28       : in  std_logic;
    l28        : out std_logic;
    l27        : out std_logic;
    ob27       : in  std_logic;
    ob26       : in  std_logic;
    l26        : out std_logic;
    l25        : out std_logic;
    ob25       : in  std_logic;
    ob24       : in  std_logic;
    lparl      : out std_logic;
    \-lparm\   : out std_logic;
    lparity    : out std_logic;
    \-lparity\ : out std_logic;
    l24        : out std_logic
    );
end;
