library ieee;
use ieee.std_logic_1164.all;

library work;
use work.other.all;

entity dip_sip180_390_8 is
  port (
    p2 : inout std_logic;
    p3 : inout std_logic;
    p4 : inout std_logic;
    p5 : inout std_logic;
    p6 : inout std_logic;
    p7 : inout std_logic
    );
end entity;

architecture dip of dip_sip180_390_8 is
begin
  -- Empty architecture as requested
end architecture;