library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ic_7437 is
  port (
    g1a : in  std_logic;
    g1b : in  std_logic;
    g1y : out std_logic;
    g2a : in  std_logic;
    g2b : in  std_logic;
    g2y : out std_logic;
    g3y : out std_logic;
    g3a : in  std_logic;
    g3b : in  std_logic;
    g4y : out std_logic;
    g4a : in  std_logic;
    g4b : in  std_logic
    );
end ic_7437;

architecture ttl of ic_7437 is
begin

end ttl;
