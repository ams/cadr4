library ieee;
use ieee.std_logic_1164.all;

entity cadr1_dbgout is
  port (
    \-select debug\ : in     std_logic;
    \dbub master\   : in     std_logic;
    \debug ack\     : in     std_logic;
    \debug in wr\   : in     std_logic;
    \debug out ack\ : in     std_logic;
    \hi 1-14\       : in     std_logic;
    \hi 15-30\      : in     std_logic;
    \ud > debug\    : in     std_logic;
    \xbus par in\   : in     std_logic;
    uba1            : in     std_logic;
    uba2            : in     std_logic;
    uba3            : in     std_logic;
    uba4            : in     std_logic;
    ubrd            : in     std_logic;
    ubwr            : in     std_logic;
    \-dbd enb\      : inout  std_logic;
    \debug active\  : inout  std_logic;
    \select debug dlyd\ : inout  std_logic;
    \select debug\  : inout  std_logic;
    dbd0            : inout  std_logic;
    dbd1            : inout  std_logic;
    dbd10           : inout  std_logic;
    dbd11           : inout  std_logic;
    dbd12           : inout  std_logic;
    dbd13           : inout  std_logic;
    dbd14           : inout  std_logic;
    dbd15           : inout  std_logic;
    dbd2            : inout  std_logic;
    dbd3            : inout  std_logic;
    dbd4            : inout  std_logic;
    dbd5            : inout  std_logic;
    dbd6            : inout  std_logic;
    dbd7            : inout  std_logic;
    dbd8            : inout  std_logic;
    dbd9            : inout  std_logic;
    udo0            : inout  std_logic;
    udo1            : inout  std_logic;
    udo10           : inout  std_logic;
    udo11           : inout  std_logic;
    udo12           : inout  std_logic;
    udo13           : inout  std_logic;
    udo14           : inout  std_logic;
    udo15           : inout  std_logic;
    udo2            : inout  std_logic;
    udo3            : inout  std_logic;
    udo4            : inout  std_logic;
    udo5            : inout  std_logic;
    udo6            : inout  std_logic;
    udo7            : inout  std_logic;
    udo8            : inout  std_logic;
    udo9            : inout  std_logic;
    \-debug > ud\   : out    std_logic;
    \-debug out req\ : out    std_logic;
    \debug in ack\  : out    std_logic;
    \debug out a0\  : out    std_logic;
    \debug out a1\  : out    std_logic;
    \debug out wr\  : out    std_logic;
    \debug ssyn\    : out    std_logic;
    \mempar to lm\  : out    std_logic;
    \spy adr1\      : out    std_logic;
    \spy adr2\      : out    std_logic;
    \spy adr3\      : out    std_logic;
    \spy adr4\      : out    std_logic
  );
end entity cadr1_dbgout;
