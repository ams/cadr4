-- CADR1_UBA
-- Generated entity from suds architecture

library ieee;
use ieee.std_logic_1164.all;

entity cadr1_uba is
  port (
    \-ub adr0\ : inout std_logic;
    \-ub adr1\ : inout std_logic;
    \-ub adr10\ : inout std_logic;
    \-ub adr11\ : inout std_logic;
    \-ub adr12\ : inout std_logic;
    \-ub adr13\ : inout std_logic;
    \-ub adr14\ : inout std_logic;
    \-ub adr15\ : inout std_logic;
    \-ub adr16\ : inout std_logic;
    \-ub adr17\ : inout std_logic;
    \-ub adr2\ : inout std_logic;
    \-ub adr3\ : inout std_logic;
    \-ub adr4\ : inout std_logic;
    \-ub adr5\ : inout std_logic;
    \-ub adr6\ : inout std_logic;
    \-ub adr7\ : inout std_logic;
    \-ub adr8\ : inout std_logic;
    \-ub adr9\ : inout std_logic;
    \-ub c1\ : inout std_logic;
    \-uba 12\ : out std_logic;
    \-uba 14\ : out std_logic;
    \-uba 15\ : out std_logic;
    \-uba 7\ : out std_logic;
    \-uba 8\ : out std_logic;
    \-uba 9\ : out std_logic;
    \-ubadrive\ : inout std_logic;
    \c1 in\ : inout std_logic;
    \c1 out\ : inout std_logic;
    uao1 : inout std_logic;
    uao10 : inout std_logic;
    uao11 : inout std_logic;
    uao12 : inout std_logic;
    uao13 : inout std_logic;
    uao14 : inout std_logic;
    uao15 : inout std_logic;
    uao16 : inout std_logic;
    uao17 : inout std_logic;
    uao2 : inout std_logic;
    uao3 : inout std_logic;
    uao4 : inout std_logic;
    uao5 : inout std_logic;
    uao6 : inout std_logic;
    uao7 : inout std_logic;
    uao8 : inout std_logic;
    uao9 : inout std_logic;
    \uba 12\ : in std_logic;
    \uba 14\ : in std_logic;
    \uba 15\ : in std_logic;
    \uba 7\ : in std_logic;
    \uba 8\ : in std_logic;
    \uba 9\ : in std_logic;
    uba0 : inout std_logic;
    uba1 : inout std_logic;
    uba10 : inout std_logic;
    uba11 : inout std_logic;
    uba12 : inout std_logic;
    uba13 : inout std_logic;
    uba14 : inout std_logic;
    uba15 : inout std_logic;
    uba16 : inout std_logic;
    uba17 : inout std_logic;
    uba2 : inout std_logic;
    uba3 : inout std_logic;
    uba4 : inout std_logic;
    uba5 : inout std_logic;
    uba6 : inout std_logic;
    uba7 : inout std_logic;
    uba8 : inout std_logic;
    uba9 : inout std_logic
  );
end entity;
