library ieee;
use ieee.std_logic_1164.all;

entity cadr1_dbgout is
  port (
    \-select debug\ : in     std_logic;
    \dbub master\   : in     std_logic;
    \debug ack\     : in     std_logic;
    \debug in wr\   : in     std_logic;
    \debug out ack\ : in     std_logic;
    \hi 1-14\       : in     std_logic;
    \hi 15-30\      : in     std_logic;
    \select debug dlyd\ : in     std_logic;
    \ud > debug\    : in     std_logic;
    \xbus par in\   : in     std_logic;
    dbd0            : in     std_logic;
    dbd1            : in     std_logic;
    dbd10           : in     std_logic;
    dbd11           : in     std_logic;
    dbd12           : in     std_logic;
    dbd13           : in     std_logic;
    dbd14           : in     std_logic;
    dbd15           : in     std_logic;
    dbd2            : in     std_logic;
    dbd3            : in     std_logic;
    dbd4            : in     std_logic;
    dbd5            : in     std_logic;
    dbd6            : in     std_logic;
    dbd7            : in     std_logic;
    dbd8            : in     std_logic;
    dbd9            : in     std_logic;
    uba1            : in     std_logic;
    uba2            : in     std_logic;
    uba3            : in     std_logic;
    uba4            : in     std_logic;
    ubrd            : in     std_logic;
    ubwr            : in     std_logic;
    udo0            : in     std_logic;
    udo1            : in     std_logic;
    udo10           : in     std_logic;
    udo11           : in     std_logic;
    udo12           : in     std_logic;
    udo13           : in     std_logic;
    udo14           : in     std_logic;
    udo15           : in     std_logic;
    udo2            : in     std_logic;
    udo3            : in     std_logic;
    udo4            : in     std_logic;
    udo5            : in     std_logic;
    udo6            : in     std_logic;
    udo7            : in     std_logic;
    udo8            : in     std_logic;
    udo9            : in     std_logic;
    \-dbd enb\      : inout  std_logic;
    \debug active\  : inout  std_logic;
    \select debug\  : inout  std_logic;
    \-debug > ud\   : out    std_logic;
    \-debug out req\ : out    std_logic;
    \debug in ack\  : out    std_logic;
    \debug out a0\  : out    std_logic;
    \debug out a1\  : out    std_logic;
    \debug out wr\  : out    std_logic;
    \debug ssyn\    : out    std_logic;
    \mempar to lm\  : out    std_logic;
    \spy adr1\      : out    std_logic;
    \spy adr2\      : out    std_logic;
    \spy adr3\      : out    std_logic;
    \spy adr4\      : out    std_logic
  );
end entity cadr1_dbgout;
