library ieee;
use ieee.std_logic_1164.all;

entity cadr_ictl is
  port (
    ramdisable      : out std_logic;
    hi1             : in  std_logic;
    \-iwriteda\     : out std_logic;
    \-promdisabled\ : out std_logic;
    idebug          : in  std_logic;
    iwriteda        : out std_logic;
    promdisabled    : in  std_logic;
    \-wp5\          : in  std_logic;
    wp5d            : out std_logic;
    wp5c            : out std_logic;
    wp5b            : out std_logic;
    wp5a            : out std_logic;
    pc0             : in  std_logic;
    \-pcb0\         : out std_logic;
    pc1             : in  std_logic;
    \-pcb1\         : out std_logic;
    pc2             : in  std_logic;
    \-pcb2\         : out std_logic;
    \-pcb3\         : out std_logic;
    pc3             : in  std_logic;
    \-pcb4\         : out std_logic;
    pc4             : in  std_logic;
    \-pcb5\         : out std_logic;
    pc5             : in  std_logic;
    \-iwea\         : out std_logic;
    \-iweb\         : out std_logic;
    \-iwei\         : out std_logic;
    \-iwej\         : out std_logic;
    pc13            : in  std_logic;
    \-pc13b\        : out std_logic;
    pc12            : in  std_logic;
    \-pc12b\        : out std_logic;
    \-iwrited\      : in  std_logic;
    iwritedd        : out std_logic;
    iwritedc        : out std_logic;
    iwritedb        : out std_logic;
    pc6             : in  std_logic;
    \-pcb6\         : out std_logic;
    pc7             : in  std_logic;
    \-pcb7\         : out std_logic;
    pc8             : in  std_logic;
    \-pcb8\         : out std_logic;
    \-pcb9\         : out std_logic;
    pc9             : in  std_logic;
    \-pcb10\        : out std_logic;
    pc10            : in  std_logic;
    \-pcb11\        : out std_logic;
    pc11            : in  std_logic;
    \-ice3a\        : out std_logic;
    \-ice2a\        : out std_logic;
    \-ice1a\        : out std_logic;
    \-ice0a\        : out std_logic;
    \-ice0b\        : out std_logic;
    \-ice1b\        : out std_logic;
    \-ice2b\        : out std_logic;
    \-ice3b\        : out std_logic;
    \-iwec\         : out std_logic;
    \-iwed\         : out std_logic;
    \-iwek\         : out std_logic;
    \-iwel\         : out std_logic;
    \-pcc0\         : out std_logic;
    \-pcc1\         : out std_logic;
    \-pcc2\         : out std_logic;
    \-pcc3\         : out std_logic;
    \-pcc4\         : out std_logic;
    \-pcc5\         : out std_logic;
    \-pcc6\         : out std_logic;
    \-pcc7\         : out std_logic;
    \-pcc8\         : out std_logic;
    \-pcc9\         : out std_logic;
    \-pcc10\        : out std_logic;
    \-pcc11\        : out std_logic;
    \-iwee\         : out std_logic;
    \-iwef\         : out std_logic;
    \-iwem\         : out std_logic;
    \-iwen\         : out std_logic;
    \-ice3c\        : out std_logic;
    \-ice2c\        : out std_logic;
    \-ice1c\        : out std_logic;
    \-ice0c\        : out std_logic;
    \-ice0d\        : out std_logic;
    \-ice1d\        : out std_logic;
    \-ice2d\        : out std_logic;
    \-ice3d\        : out std_logic;
    \-iweg\         : out std_logic;
    \-iweh\         : out std_logic;
    \-iweo\         : out std_logic;
    \-iwep\         : out std_logic);
end;
