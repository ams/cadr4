library ieee;
use ieee.std_logic_1164.all;

entity cadr_pdl0 is
  port (
    \-pdla0b\       : in     std_logic;
    \-pdla1b\       : in     std_logic;
    \-pdla2b\       : in     std_logic;
    \-pdla3b\       : in     std_logic;
    \-pdla4b\       : in     std_logic;
    \-pdla5b\       : in     std_logic;
    \-pdla6b\       : in     std_logic;
    \-pdla7b\       : in     std_logic;
    \-pdla8b\       : in     std_logic;
    \-pdla9b\       : in     std_logic;
    \-pwpa\         : in     std_logic;
    \-pwpb\         : in     std_logic;
    l16             : in     std_logic;
    l17             : in     std_logic;
    l18             : in     std_logic;
    l19             : in     std_logic;
    l20             : in     std_logic;
    l21             : in     std_logic;
    l22             : in     std_logic;
    l23             : in     std_logic;
    l24             : in     std_logic;
    l25             : in     std_logic;
    l26             : in     std_logic;
    l27             : in     std_logic;
    l28             : in     std_logic;
    l29             : in     std_logic;
    l30             : in     std_logic;
    l31             : in     std_logic;
    lparity         : in     std_logic;
    pdl16           : out    std_logic;
    pdl17           : out    std_logic;
    pdl18           : out    std_logic;
    pdl19           : out    std_logic;
    pdl20           : out    std_logic;
    pdl21           : out    std_logic;
    pdl22           : out    std_logic;
    pdl23           : out    std_logic;
    pdl24           : out    std_logic;
    pdl25           : out    std_logic;
    pdl26           : out    std_logic;
    pdl27           : out    std_logic;
    pdl28           : out    std_logic;
    pdl29           : out    std_logic;
    pdl30           : out    std_logic;
    pdl31           : out    std_logic;
    pdlparity       : out    std_logic
  );
end entity cadr_pdl0;
