library ieee;
use ieee.std_logic_1164.all;

entity helper_deassert_halt is
  port (
    \-halt\: out std_logic := '1'
  );
end entity;

architecture structural of helper_deassert_halt is
begin
end architecture;