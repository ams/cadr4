library ieee;
use ieee.std_logic_1164.all;

entity busint_ubmap is
  port (
    \-ubmap > udo\  : in     std_logic;
    \-ubmapwe\      : in     std_logic;
    \select page\   : in     std_logic;
    uba1            : in     std_logic;
    uba10           : in     std_logic;
    uba11           : in     std_logic;
    uba12           : in     std_logic;
    uba13           : in     std_logic;
    uba2            : in     std_logic;
    uba3            : in     std_logic;
    uba4            : in     std_logic;
    udi0            : in     std_logic;
    udi1            : in     std_logic;
    udi10           : in     std_logic;
    udi11           : in     std_logic;
    udi12           : in     std_logic;
    udi13           : in     std_logic;
    udi14           : in     std_logic;
    udi15           : in     std_logic;
    udi2            : in     std_logic;
    udi3            : in     std_logic;
    udi4            : in     std_logic;
    udi5            : in     std_logic;
    udi6            : in     std_logic;
    udi7            : in     std_logic;
    udi8            : in     std_logic;
    udi9            : in     std_logic;
    \-ubpn0a\       : out    std_logic;
    \-ubpn0b\       : out    std_logic;
    \-ubpn1a\       : out    std_logic;
    \-ubpn1b\       : out    std_logic;
    \-ubpn2a\       : out    std_logic;
    \-ubpn2b\       : out    std_logic;
    \-ubpn3a\       : out    std_logic;
    \-ubpn3b\       : out    std_logic;
    mapvalid        : out    std_logic;
    ubma10          : out    std_logic;
    ubma11          : out    std_logic;
    ubma12          : out    std_logic;
    ubma13          : out    std_logic;
    ubma14          : out    std_logic;
    ubma15          : out    std_logic;
    ubma16          : out    std_logic;
    ubma17          : out    std_logic;
    ubma18          : out    std_logic;
    ubma19          : out    std_logic;
    ubma20          : out    std_logic;
    ubma21          : out    std_logic;
    ubma8           : out    std_logic;
    ubma9           : out    std_logic;
    udo0            : out    std_logic;
    udo1            : out    std_logic;
    udo10           : out    std_logic;
    udo11           : out    std_logic;
    udo12           : out    std_logic;
    udo13           : out    std_logic;
    udo14           : out    std_logic;
    udo15           : out    std_logic;
    udo2            : out    std_logic;
    udo3            : out    std_logic;
    udo4            : out    std_logic;
    udo5            : out    std_logic;
    udo6            : out    std_logic;
    udo7            : out    std_logic;
    udo8            : out    std_logic;
    udo9            : out    std_logic;
    writeok         : out    std_logic
  );
end entity;
