library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_qctl is
  port (
    \-qdrive\ : out std_logic;
    tse2      : in  std_logic;
    srcq      : out std_logic;
    q7        : in  std_logic;
    mf0       : out std_logic;
    q6        : in  std_logic;
    mf1       : out std_logic;
    q5        : in  std_logic;
    mf2       : out std_logic;
    q4        : in  std_logic;
    mf3       : out std_logic;
    q3        : in  std_logic;
    mf4       : out std_logic;
    q2        : in  std_logic;
    mf5       : out std_logic;
    q1        : in  std_logic;
    mf6       : out std_logic;
    q0        : in  std_logic;
    mf7       : out std_logic;
    qdrive    : out std_logic;
    q31       : in  std_logic;
    mf24      : out std_logic;
    q30       : in  std_logic;
    mf25      : out std_logic;
    q29       : in  std_logic;
    mf26      : out std_logic;
    q28       : in  std_logic;
    mf27      : out std_logic;
    q27       : in  std_logic;
    mf28      : out std_logic;
    q26       : in  std_logic;
    mf29      : out std_logic;
    q25       : in  std_logic;
    mf30      : out std_logic;
    q24       : in  std_logic;
    mf31      : out std_logic;
    q23       : in  std_logic;
    mf16      : out std_logic;
    q22       : in  std_logic;
    mf17      : out std_logic;
    q21       : in  std_logic;
    mf18      : out std_logic;
    q20       : in  std_logic;
    mf19      : out std_logic;
    q19       : in  std_logic;
    mf20      : out std_logic;
    q18       : in  std_logic;
    mf21      : out std_logic;
    q17       : in  std_logic;
    mf22      : out std_logic;
    q16       : in  std_logic;
    mf23      : out std_logic;
    q15       : in  std_logic;
    mf8       : out std_logic;
    q14       : in  std_logic;
    mf9       : out std_logic;
    q13       : in  std_logic;
    mf10      : out std_logic;
    q12       : in  std_logic;
    mf11      : out std_logic;
    q11       : in  std_logic;
    mf12      : out std_logic;
    q10       : in  std_logic;
    mf13      : out std_logic;
    q9        : in  std_logic;
    mf14      : out std_logic;
    q8        : in  std_logic;
    mf15      : out std_logic;
    \-srcq\   : in  std_logic;
    \-alu31\  : out std_logic;
    alu31     : in  std_logic;
    \-iralu\  : in  std_logic;
    \-ir1\    : in  std_logic;
    qs1       : out std_logic;
    \-ir0\    : in  std_logic;
    qs0       : out std_logic);
end;

architecture ttl of cadr_qctl is
begin
  qctl_1a18 : sn74s00 port map(g3q_n   => \-qdrive\, g3b => tse2, g3a => srcq, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g4a => '0', g4b => '0');
  qctl_1e12 : sn74s241 port map(aenb_n => \-qdrive\, ain0 => q7, bout3 => mf0, ain1 => q6, bout2 => mf1, ain2 => q5, bout1 => mf2, ain3 => q4, bout0 => mf3, bin0 => q3, aout3 => mf4, bin1 => q2, aout2 => mf5, bin2 => q1, aout1 => mf6, bin3 => q0, aout0 => mf7, benb => qdrive);
  qctl_1f08 : sn74s241 port map(aenb_n => \-qdrive\, ain0 => q31, bout3 => mf24, ain1 => q30, bout2 => mf25, ain2 => q29, bout1 => mf26, ain3 => q28, bout0 => mf27, bin0 => q27, aout3 => mf28, bin1 => q26, aout2 => mf29, bin2 => q25, aout1 => mf30, bin3 => q24, aout0 => mf31, benb => qdrive);
  qctl_1f10 : sn74s241 port map(aenb_n => \-qdrive\, ain0 => q23, bout3 => mf16, ain1 => q22, bout2 => mf17, ain2 => q21, bout1 => mf18, ain3 => q20, bout0 => mf19, bin0 => q19, aout3 => mf20, bin1 => q18, aout2 => mf21, bin2 => q17, aout1 => mf22, bin3 => q16, aout0 => mf23, benb => qdrive);
  qctl_1f15 : sn74s241 port map(aenb_n => \-qdrive\, ain0 => q15, bout3 => mf8, ain1 => q14, bout2 => mf9, ain2 => q13, bout1 => mf10, ain3 => q12, bout0 => mf11, bin0 => q11, aout3 => mf12, bin1 => q10, aout2 => mf13, bin2 => q9, aout1 => mf14, bin3 => q8, aout0 => mf15, benb => qdrive);
  qctl_2a04 : sn74s08 port map(g4q     => qdrive, g4a => tse2, g4b => srcq, g1b => '0', g1a => '0', g2b => '0', g2a => '0', g3a => '0', g3b => '0');
  qctl_2a05 : sn74s04 port map(g5q_n   => srcq, g5a => \-srcq\, g6q_n => \-alu31\, g6a => alu31, g1a => '0', g2a => '0', g3a => '0', g4a => '0');
  qctl_2b19 : sn7428 port map(g3a      => \-iralu\, g3b => \-ir1\, g3q_n => qs1, g4a => \-iralu\, g4b => \-ir0\, g4q_n => qs0, g1a => '0', g1b => '0', g2a => '0', g2b => '0');
end architecture;
