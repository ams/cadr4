library ieee;
use ieee.std_logic_1164.all;

entity cadr1_lmdata is
  port (
    \-lmbus enb\    : in     std_logic;
    \bus > lm\      : in     std_logic;
    bus0            : inout  std_logic;
    bus1            : inout  std_logic;
    bus10           : inout  std_logic;
    bus11           : inout  std_logic;
    bus12           : inout  std_logic;
    bus13           : inout  std_logic;
    bus14           : inout  std_logic;
    bus15           : inout  std_logic;
    bus16           : inout  std_logic;
    bus17           : inout  std_logic;
    bus18           : inout  std_logic;
    bus19           : inout  std_logic;
    bus2            : inout  std_logic;
    bus20           : inout  std_logic;
    bus21           : inout  std_logic;
    bus22           : inout  std_logic;
    bus23           : inout  std_logic;
    bus24           : inout  std_logic;
    bus25           : inout  std_logic;
    bus26           : inout  std_logic;
    bus27           : inout  std_logic;
    bus28           : inout  std_logic;
    bus29           : inout  std_logic;
    bus3            : inout  std_logic;
    bus30           : inout  std_logic;
    bus31           : inout  std_logic;
    bus4            : inout  std_logic;
    bus5            : inout  std_logic;
    bus6            : inout  std_logic;
    bus7            : inout  std_logic;
    bus8            : inout  std_logic;
    bus9            : inout  std_logic;
    mem0            : inout  std_logic;
    mem1            : inout  std_logic;
    mem10           : inout  std_logic;
    mem11           : inout  std_logic;
    mem12           : inout  std_logic;
    mem13           : inout  std_logic;
    mem14           : inout  std_logic;
    mem15           : inout  std_logic;
    mem16           : inout  std_logic;
    mem17           : inout  std_logic;
    mem18           : inout  std_logic;
    mem19           : inout  std_logic;
    mem2            : inout  std_logic;
    mem20           : inout  std_logic;
    mem21           : inout  std_logic;
    mem22           : inout  std_logic;
    mem23           : inout  std_logic;
    mem24           : inout  std_logic;
    mem25           : inout  std_logic;
    mem26           : inout  std_logic;
    mem27           : inout  std_logic;
    mem28           : inout  std_logic;
    mem29           : inout  std_logic;
    mem3            : inout  std_logic;
    mem30           : inout  std_logic;
    mem31           : inout  std_logic;
    mem4            : inout  std_logic;
    mem5            : inout  std_logic;
    mem6            : inout  std_logic;
    mem7            : inout  std_logic;
    mem8            : inout  std_logic;
    mem9            : inout  std_logic
  );
end entity cadr1_lmdata;
