library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity res20 is
  port (
    r2  : out std_logic;
    r3  : out std_logic;
    r4  : out std_logic;
    r5  : out std_logic;
    r6  : out std_logic;
    r7  : out std_logic;
    r8  : out std_logic;
    r9  : out std_logic;
    r10 : out std_logic;
    r11 : out std_logic;
    r12 : out std_logic;
    r13 : out std_logic;
    r14 : out std_logic;
    r15 : out std_logic;
    r16 : out std_logic;
    r17 : out std_logic;
    r18 : out std_logic;
    r19 : out std_logic
    );
end;

-- ChatGPT Codex implementation
architecture ttl of res20 is
begin
  r2  <= '1'; r3  <= '1'; r4  <= '1'; r5  <= '1';
  r6  <= '1'; r7  <= '1'; r8  <= '1'; r9  <= '1';
  r10 <= '1'; r11 <= '1'; r12 <= '1'; r13 <= '1';
  r14 <= '1'; r15 <= '1'; r16 <= '1'; r17 <= '1';
  r18 <= '1'; r19 <= '1';
end;
