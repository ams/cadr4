library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.sn74.all;

entity sn74181_tb is
end;

architecture testbench of sn74181_tb is

  -- Initialize signals to avoid metavalue assertions
  signal cin_n  : std_logic := '1';
  signal s0     : std_logic := '0';
  signal s1     : std_logic := '0';
  signal s2     : std_logic := '0';
  signal s3     : std_logic := '0';
  signal m      : std_logic := '0';
  signal a0     : std_logic := '0';
  signal a1     : std_logic := '0';
  signal a2     : std_logic := '0';
  signal a3     : std_logic := '0';
  signal b0     : std_logic := '0';
  signal b1     : std_logic := '0';
  signal b2     : std_logic := '0';
  signal b3     : std_logic := '0';
  signal f0     : std_logic;
  signal f1     : std_logic;
  signal f2     : std_logic;
  signal f3     : std_logic;
  signal aeb    : std_logic;
  signal x      : std_logic;
  signal y      : std_logic;
  signal cout_n : std_logic;

begin

  uut : sn74181 port map(
    cout_n => cout_n,
    y      => y,
    x      => x,
    aeb    => aeb,
    f3     => f3,
    f2     => f2,
    f1     => f1,
    f0     => f0,
    b3     => b3,
    b2     => b2,
    b1     => b1,
    b0     => b0,
    a3     => a3,
    a2     => a2,
    a1     => a1,
    a0     => a0,
    m      => m,
    s3     => s3,
    s2     => s2,
    s1     => s1,
    s0     => s0,
    cin_n  => cin_n
  );

  process
    variable f_result : std_logic_vector(3 downto 0);
  begin
    
    -- Test Logic Mode (M = 1) - Table 2 Active High Data
    report "Testing Logic Mode (M=1)";
    m <= '1';
    cin_n <= '1'; -- Don't care in logic mode
    
    -- Test data: A=1010 (10), B=0110 (6)
    a3 <= '1'; a2 <= '0'; a1 <= '1'; a0 <= '0'; -- A=10
    b3 <= '0'; b2 <= '1'; b1 <= '1'; b0 <= '0'; -- B=6
    
    -- S=0000: F = NOT A
    s3 <= '0'; s2 <= '0'; s1 <= '0'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0101" report "Logic S=0000 (NOT A) failed" severity error;
    
    -- S=0001: F = NOT(A+B)
    s3 <= '0'; s2 <= '0'; s1 <= '0'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0001" report "Logic S=0001 (NOT(A+B)) failed" severity error;
    
    -- S=0010: F = (NOT A)B
    s3 <= '0'; s2 <= '0'; s1 <= '1'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0100" report "Logic S=0010 ((NOT A)B) failed" severity error;
    
    -- S=0011: F = 0
    s3 <= '0'; s2 <= '0'; s1 <= '1'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0000" report "Logic S=0011 (0) failed" severity error;
    
    -- S=0100: F = NOT(AB)
    s3 <= '0'; s2 <= '1'; s1 <= '0'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1101" report "Logic S=0100 (NOT(AB)) failed" severity error;
    
    -- S=0101: F = NOT B
    s3 <= '0'; s2 <= '1'; s1 <= '0'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1001" report "Logic S=0101 (NOT B) failed" severity error;
    
    -- S=0110: F = A XOR B
    s3 <= '0'; s2 <= '1'; s1 <= '1'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1100" report "Logic S=0110 (A XOR B) failed" severity error;
    
    -- S=0111: F = A(NOT B)
    s3 <= '0'; s2 <= '1'; s1 <= '1'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1000" report "Logic S=0111 (A(NOT B)) failed" severity error;
    
    -- S=1000: F = (NOT A)+B
    s3 <= '1'; s2 <= '0'; s1 <= '0'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0111" report "Logic S=1000 ((NOT A)+B) failed" severity error;
    
    -- S=1001: F = NOT(A XOR B)
    s3 <= '1'; s2 <= '0'; s1 <= '0'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0011" report "Logic S=1001 (NOT(A XOR B)) failed" severity error;
    
    -- S=1010: F = B
    s3 <= '1'; s2 <= '0'; s1 <= '1'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0110" report "Logic S=1010 (B) failed" severity error;
    
    -- S=1011: F = AB
    s3 <= '1'; s2 <= '0'; s1 <= '1'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0010" report "Logic S=1011 (AB) failed" severity error;
    
    -- S=1100: F = 1
    s3 <= '1'; s2 <= '1'; s1 <= '0'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1111" report "Logic S=1100 (1) failed" severity error;
    
    -- S=1101: F = A+(NOT B)
    s3 <= '1'; s2 <= '1'; s1 <= '0'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1011" report "Logic S=1101 (A+(NOT B)) failed" severity error;
    
    -- S=1110: F = A+B
    s3 <= '1'; s2 <= '1'; s1 <= '1'; s0 <= '0';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1110" report "Logic S=1110 (A+B) failed" severity error;
    
    -- S=1111: F = A
    s3 <= '1'; s2 <= '1'; s1 <= '1'; s0 <= '1';
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1010" report "Logic S=1111 (A) failed" severity error;
    
    -- Test Arithmetic Mode (M = 0) - Table 2 Active High Data
    report "Testing Arithmetic Mode (M=0)";
    m <= '0';
    
    -- Test data: A=5 (0101), B=3 (0011)
    a3 <= '0'; a2 <= '1'; a1 <= '0'; a0 <= '1'; -- A=5
    b3 <= '0'; b2 <= '0'; b1 <= '1'; b0 <= '1'; -- B=3
    
    -- S=0000: F = A (Cn=0) / A+1 (Cn=1)
    s3 <= '0'; s2 <= '0'; s1 <= '0'; s0 <= '0';
    cin_n <= '1'; -- Cn=0
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0101" report "Arith S=0000 Cn=0 (A) failed" severity error;
    
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0110" report "Arith S=0000 Cn=1 (A+1) failed" severity error;
    
    -- S=0001: F = A+B (Cn=0) / A+B+1 (Cn=1)
    s3 <= '0'; s2 <= '0'; s1 <= '0'; s0 <= '1';
    cin_n <= '1'; -- Cn=0
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1000" report "Arith S=0001 Cn=0 (A+B) failed" severity error;
    
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1001" report "Arith S=0001 Cn=1 (A+B+1) failed" severity error;
    
    -- S=0010: F = A+(NOT B) (Cn=0) / A+(NOT B)+1 (Cn=1)
    s3 <= '0'; s2 <= '0'; s1 <= '1'; s0 <= '0';
    cin_n <= '1'; -- Cn=0
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0001" report "Arith S=0010 Cn=0 (A+(NOT B)) failed" severity error;
    
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0010" report "Arith S=0010 Cn=1 (A-B) failed" severity error;
    
    -- S=0110: F = A-B-1 (Cn=0) / A-B (Cn=1)
    s3 <= '0'; s2 <= '1'; s1 <= '1'; s0 <= '0';
    cin_n <= '1'; -- Cn=0
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0001" report "Arith S=0110 Cn=0 (A-B-1) failed" severity error;
    
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0010" report "Arith S=0110 Cn=1 (A-B) failed" severity error;
    
    -- S=1100: F = A+A (Cn=0) / A+A+1 (Cn=1) [shift left]
    s3 <= '1'; s2 <= '1'; s1 <= '0'; s0 <= '0';
    cin_n <= '1'; -- Cn=0
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1010" report "Arith S=1100 Cn=0 (A+A) failed" severity error;
    
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "1011" report "Arith S=1100 Cn=1 (A+A+1) failed" severity error;
    
    -- S=1111: F = A-1 (Cn=0) / A (Cn=1)
    s3 <= '1'; s2 <= '1'; s1 <= '1'; s0 <= '1';
    cin_n <= '1'; -- Cn=0
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0100" report "Arith S=1111 Cn=0 (A-1) failed" severity error;
    
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    f_result := f3 & f2 & f1 & f0;
    assert f_result = "0101" report "Arith S=1111 Cn=1 (A) failed" severity error;
    
    -- Test A equals B
    report "Testing A equals B";
    a3 <= '0'; a2 <= '1'; a1 <= '0'; a0 <= '1'; -- A=5
    b3 <= '0'; b2 <= '1'; b1 <= '0'; b0 <= '1'; -- B=5
    wait for 10 ns;
    assert aeb = '1' report "A equals B failed when A=B=5" severity error;
    
    a3 <= '0'; a2 <= '1'; a1 <= '0'; a0 <= '1'; -- A=5
    b3 <= '0'; b2 <= '0'; b1 <= '1'; b0 <= '1'; -- B=3
    wait for 10 ns;
    assert aeb = '0' report "A equals B failed when A=5, B=3" severity error;
    
    -- Test carry propagate (X) and carry generate (Y)
    report "Testing carry propagate and generate";
    m <= '0'; -- Arithmetic mode
    a3 <= '1'; a2 <= '1'; a1 <= '1'; a0 <= '1'; -- A=15
    b3 <= '0'; b2 <= '0'; b1 <= '0'; b0 <= '1'; -- B=1
    s3 <= '0'; s2 <= '0'; s1 <= '0'; s0 <= '1'; -- A+B
    cin_n <= '0'; -- Cn=1
    wait for 10 ns;
    -- This should generate carry out (Y=1) and overflow
    assert cout_n = '0' report "Carry out should be active (cout_n=0) for 15+1+1" severity error;
    
    report "All tests completed successfully";
    wait;
  end process;

end;
