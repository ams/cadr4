library ieee;
use ieee.std_logic_1164.all;

entity cadr_mf is
  port (
    tse1a      : in  std_logic;
    mfenb      : out std_logic;
    \-mfdrive\ : out std_logic;
    mf23       : in  std_logic;
    m16        : out std_logic;
    mf22       : in  std_logic;
    m17        : out std_logic;
    mf21       : in  std_logic;
    m18        : out std_logic;
    mf20       : in  std_logic;
    m19        : out std_logic;
    mf19       : in  std_logic;
    m20        : out std_logic;
    mf18       : in  std_logic;
    m21        : out std_logic;
    mf17       : in  std_logic;
    m22        : out std_logic;
    mf16       : in  std_logic;
    m23        : out std_logic;
    mfdrive    : out std_logic;
    mf15       : in  std_logic;
    m8         : out std_logic;
    mf14       : in  std_logic;
    m9         : out std_logic;
    mf13       : in  std_logic;
    m10        : out std_logic;
    mf12       : in  std_logic;
    m11        : out std_logic;
    mf11       : in  std_logic;
    m12        : out std_logic;
    mf10       : in  std_logic;
    m13        : out std_logic;
    mf9        : in  std_logic;
    m14        : out std_logic;
    mf8        : in  std_logic;
    m15        : out std_logic;
    mf7        : in  std_logic;
    m0         : out std_logic;
    mf6        : in  std_logic;
    m1         : out std_logic;
    mf5        : in  std_logic;
    m2         : out std_logic;
    mf4        : in  std_logic;
    m3         : out std_logic;
    mf3        : in  std_logic;
    m4         : out std_logic;
    mf2        : in  std_logic;
    m5         : out std_logic;
    mf1        : in  std_logic;
    m6         : out std_logic;
    mf0        : in  std_logic;
    m7         : out std_logic;
    mf31       : in  std_logic;
    m24        : out std_logic;
    mf30       : in  std_logic;
    m25        : out std_logic;
    mf29       : in  std_logic;
    m26        : out std_logic;
    mf28       : in  std_logic;
    m27        : out std_logic;
    mf27       : in  std_logic;
    m28        : out std_logic;
    mf26       : in  std_logic;
    m29        : out std_logic;
    mf25       : in  std_logic;
    m30        : out std_logic;
    mf24       : in  std_logic;
    m31        : out std_logic;
    pdlenb     : in  std_logic;
    spcenb     : in  std_logic;
    \-srcm\    : out std_logic;
    \-ir31\    : in  std_logic;
    \-mpass\   : in  std_logic
    );
end;
