library ieee;
use ieee.std_logic_1164.all;

entity cadr1_dbgin is
  port (
    \-dbub master\  : in     std_logic;
    \-lm power reset\ : in     std_logic;
    \-lm unibus reset\ : in     std_logic;
    \dbub master\   : in     std_logic;
    \hi 1-14\       : in     std_logic;
    \hi 15-30\      : in     std_logic;
    \ssyn t0\       : in     std_logic;
    \unibus init in\ : in     std_logic;
    dbd0            : in     std_logic;
    dbd1            : in     std_logic;
    dbd10           : in     std_logic;
    dbd11           : in     std_logic;
    dbd12           : in     std_logic;
    dbd13           : in     std_logic;
    dbd14           : in     std_logic;
    dbd15           : in     std_logic;
    dbd2            : in     std_logic;
    dbd3            : in     std_logic;
    dbd4            : in     std_logic;
    dbd5            : in     std_logic;
    dbd6            : in     std_logic;
    dbd7            : in     std_logic;
    dbd8            : in     std_logic;
    dbd9            : in     std_logic;
    \-db adr0 clk\  : inout  std_logic;
    \-db adr1 clk\  : inout  std_logic;
    \-db need ub\   : inout  std_logic;
    \-db read status\ : inout  std_logic;
    \-debug in req\ : inout  std_logic;
    \-debug reset\  : inout  std_logic;
    \-debugee reset\ : inout  std_logic;
    \-local enable\ : inout  std_logic;
    \debug in a0\   : inout  std_logic;
    \debug in a1\   : inout  std_logic;
    \debug in wr\   : inout  std_logic;
    \debug out ack\ : inout  std_logic;
    \local enable\  : inout  std_logic;
    reset           : inout  std_logic;
    \-busint lm reset\ : out    std_logic;
    \-debug timeout inh\ : out    std_logic;
    \-reset\        : out    std_logic;
    \db need ub\    : out    std_logic;
    \debug ack\     : out    std_logic;
    uao1            : out    std_logic;
    uao10           : out    std_logic;
    uao11           : out    std_logic;
    uao12           : out    std_logic;
    uao13           : out    std_logic;
    uao14           : out    std_logic;
    uao15           : out    std_logic;
    uao16           : out    std_logic;
    uao17           : out    std_logic;
    uao2            : out    std_logic;
    uao3            : out    std_logic;
    uao4            : out    std_logic;
    uao5            : out    std_logic;
    uao6            : out    std_logic;
    uao7            : out    std_logic;
    uao8            : out    std_logic;
    uao9            : out    std_logic
  );
end entity cadr1_dbgin;
