library ieee;
use ieee.std_logic_1164.all;

use work.set.all;

entity set_tb is
end entity;

architecture structural of set_tb is
  signal \-ape\: std_logic;
  signal \-clk2c\: std_logic;
  signal \-clk3g\: std_logic;
  signal \-clk4e\: std_logic;
  signal \-clk5\: std_logic;
  signal \-clock reset b\: std_logic;
  signal \-destimod0\: std_logic;
  signal \-destimod1\: std_logic;
  signal \-destintctl\: std_logic;
  signal \-destlc\: std_logic;
  signal \-destmdr\: std_logic;
  signal \-destmem\: std_logic;
  signal \-destpdl(p)\: std_logic;
  signal \-destpdl(x)\: std_logic;
  signal \-destpdlp\: std_logic;
  signal \-destpdltop\: std_logic;
  signal \-destpdlx\: std_logic;
  signal \-destspc\: std_logic;
  signal \-destvma\: std_logic;
  signal \-div\: std_logic;
  signal \-dpe\: std_logic;
  signal \-funct2\: std_logic;
  signal \-hang\: std_logic;
  signal \-higherr\: std_logic;
  signal \-idebug\: std_logic;
  signal \-ifetch\: std_logic;
  signal \-ilong\: std_logic;
  signal \-ipe\: std_logic;
  signal \-ir0\: std_logic;
  signal \-ir12\: std_logic;
  signal \-ir13\: std_logic;
  signal \-ir1\: std_logic;
  signal \-ir2\: std_logic;
  signal \-ir31\: std_logic;
  signal \-ir3\: std_logic;
  signal \-ir4\: std_logic;
  signal \-iralu\: std_logic;
  signal \-irbyte\: std_logic;
  signal \-irdisp\: std_logic;
  signal \-irjump\: std_logic;
  signal \-iwrited\: std_logic;
  signal \-iwriteda\: std_logic;
  signal \-jcond\: std_logic;
  signal \-lcry3\: std_logic;
  signal \-ldclk\: std_logic;
  signal \-lddbirh\: std_logic;
  signal \-lddbirl\: std_logic;
  signal \-lddbirm\: std_logic;
  signal \-ldmode\: std_logic;
  signal \-ldopc\: std_logic;
  signal \-ldstat\: std_logic;
  signal \-lvmo22\: std_logic;
  signal \-lvmo23\: std_logic;
  signal \-machruna\: std_logic;
  signal \-md0\: std_logic;
  signal \-md10\: std_logic;
  signal \-md11\: std_logic;
  signal \-md12\: std_logic;
  signal \-md13\: std_logic;
  signal \-md14\: std_logic;
  signal \-md15\: std_logic;
  signal \-md16\: std_logic;
  signal \-md17\: std_logic;
  signal \-md18\: std_logic;
  signal \-md19\: std_logic;
  signal \-md1\: std_logic;
  signal \-md20\: std_logic;
  signal \-md21\: std_logic;
  signal \-md22\: std_logic;
  signal \-md23\: std_logic;
  signal \-md24\: std_logic;
  signal \-md25\: std_logic;
  signal \-md26\: std_logic;
  signal \-md27\: std_logic;
  signal \-md28\: std_logic;
  signal \-md29\: std_logic;
  signal \-md2\: std_logic;
  signal \-md30\: std_logic;
  signal \-md31\: std_logic;
  signal \-md3\: std_logic;
  signal \-md4\: std_logic;
  signal \-md5\: std_logic;
  signal \-md6\: std_logic;
  signal \-md7\: std_logic;
  signal \-md8\: std_logic;
  signal \-md9\: std_logic;
  signal \-memdrive.a\: std_logic;
  signal \-memdrive.b\: std_logic;
  signal \-mempe\: std_logic;
  signal \-memstart\: std_logic;
  signal \-mpe\: std_logic;
  signal \-mul\: std_logic;
  signal \-nop11\: std_logic;
  signal \-nopa\: std_logic;
  signal \-opcinh\: std_logic;
  signal \-pdlpe\: std_logic;
  signal \-pfr\: std_logic;
  signal \-pfw\: std_logic;
  signal \-promdisabled\: std_logic;
  signal \-reset\: std_logic;
  signal \-sh3\: std_logic;
  signal \-sh4\: std_logic;
  signal \-spcdrive\: std_logic;
  signal \-spcnt\: std_logic;
  signal \-spcpass\: std_logic;
  signal \-spcwpass\: std_logic;
  signal \-spe\: std_logic;
  signal \-spop\: std_logic;
  signal \-spy.sth\: std_logic;
  signal \-spy.stl\: std_logic;
  signal \-srcdc\: std_logic;
  signal \-srclc\: std_logic;
  signal \-srcmap\: std_logic;
  signal \-srcmd\: std_logic;
  signal \-srcopc\: std_logic;
  signal \-srcpdlidx\: std_logic;
  signal \-srcpdlpop\: std_logic;
  signal \-srcpdlptr\: std_logic;
  signal \-srcpdltop\: std_logic;
  signal \-srcq\: std_logic;
  signal \-srcspc\: std_logic;
  signal \-srcspcpop\: std_logic;
  signal \-srcspcpopreal\: std_logic;
  signal \-srcvma\: std_logic;
  signal \-statbit\: std_logic;
  signal \-stathalt\: std_logic;
  signal \-stc32\: std_logic;
  signal \-swpa\: std_logic;
  signal \-swpb\: std_logic;
  signal \-tpr60\: std_logic;
  signal \-trap\: std_logic;
  signal \-upperhighok\: std_logic;
  signal \-v0pe\: std_logic;
  signal \-v1pe\: std_logic;
  signal \-vm0wpa\: std_logic;
  signal \-vm0wpb\: std_logic;
  signal \-vm1wpa\: std_logic;
  signal \-vm1wpb\: std_logic;
  signal \-vma0\: std_logic;
  signal \-vma10\: std_logic;
  signal \-vma11\: std_logic;
  signal \-vma12\: std_logic;
  signal \-vma13\: std_logic;
  signal \-vma14\: std_logic;
  signal \-vma15\: std_logic;
  signal \-vma16\: std_logic;
  signal \-vma17\: std_logic;
  signal \-vma18\: std_logic;
  signal \-vma19\: std_logic;
  signal \-vma1\: std_logic;
  signal \-vma20\: std_logic;
  signal \-vma21\: std_logic;
  signal \-vma22\: std_logic;
  signal \-vma23\: std_logic;
  signal \-vma25\: std_logic;
  signal \-vma26\: std_logic;
  signal \-vma27\: std_logic;
  signal \-vma28\: std_logic;
  signal \-vma29\: std_logic;
  signal \-vma2\: std_logic;
  signal \-vma30\: std_logic;
  signal \-vma31\: std_logic;
  signal \-vma3\: std_logic;
  signal \-vma4\: std_logic;
  signal \-vma5\: std_logic;
  signal \-vma6\: std_logic;
  signal \-vma7\: std_logic;
  signal \-vma8\: std_logic;
  signal \-vma9\: std_logic;
  signal \-vmaenb\: std_logic;
  signal \-vmaok\: std_logic;
  signal \-vmo18\: std_logic;
  signal \-vmo19\: std_logic;
  signal \-wait\: std_logic;
  signal \-wp5\: std_logic;
  signal \a=m\: std_logic;
  signal \boot.trap\: std_logic;
  signal \int.enable\: std_logic;
  signal \lc byte mode\: std_logic;
  signal \lpc.hold\: std_logic;
  signal \prog.unibus.reset\: std_logic;
  signal \sequence.break\: std_logic;
  signal \use.md\: std_logic;
  signal a0: std_logic;
  signal a10: std_logic;
  signal a11: std_logic;
  signal a12: std_logic;
  signal a13: std_logic;
  signal a14: std_logic;
  signal a15: std_logic;
  signal a16: std_logic;
  signal a17: std_logic;
  signal a18: std_logic;
  signal a19: std_logic;
  signal a1: std_logic;
  signal a20: std_logic;
  signal a21: std_logic;
  signal a22: std_logic;
  signal a23: std_logic;
  signal a24: std_logic;
  signal a25: std_logic;
  signal a26: std_logic;
  signal a27: std_logic;
  signal a28: std_logic;
  signal a29: std_logic;
  signal a2: std_logic;
  signal a30: std_logic;
  signal a31a: std_logic;
  signal a31b: std_logic;
  signal a3: std_logic;
  signal a4: std_logic;
  signal a5: std_logic;
  signal a6: std_logic;
  signal a7: std_logic;
  signal a8: std_logic;
  signal a9: std_logic;
  signal aa0: std_logic;
  signal aa10: std_logic;
  signal aa11: std_logic;
  signal aa12: std_logic;
  signal aa13: std_logic;
  signal aa14: std_logic;
  signal aa15: std_logic;
  signal aa1: std_logic;
  signal aa2: std_logic;
  signal aa3: std_logic;
  signal aa4: std_logic;
  signal aa5: std_logic;
  signal aa6: std_logic;
  signal aa7: std_logic;
  signal aa8: std_logic;
  signal aa9: std_logic;
  signal alu0: std_logic;
  signal alu10: std_logic;
  signal alu11: std_logic;
  signal alu12: std_logic;
  signal alu13: std_logic;
  signal alu14: std_logic;
  signal alu15: std_logic;
  signal alu16: std_logic;
  signal alu17: std_logic;
  signal alu18: std_logic;
  signal alu19: std_logic;
  signal alu1: std_logic;
  signal alu20: std_logic;
  signal alu21: std_logic;
  signal alu22: std_logic;
  signal alu23: std_logic;
  signal alu24: std_logic;
  signal alu25: std_logic;
  signal alu26: std_logic;
  signal alu27: std_logic;
  signal alu28: std_logic;
  signal alu29: std_logic;
  signal alu2: std_logic;
  signal alu30: std_logic;
  signal alu31: std_logic;
  signal alu32: std_logic;
  signal alu3: std_logic;
  signal alu4: std_logic;
  signal alu5: std_logic;
  signal alu6: std_logic;
  signal alu7: std_logic;
  signal alu8: std_logic;
  signal alu9: std_logic;
  signal aparity: std_logic;
  signal aparok: std_logic;
  signal clk1a: std_logic;
  signal clk2a: std_logic;
  signal clk2b: std_logic;
  signal clk2c: std_logic;
  signal clk3a: std_logic;
  signal clk3b: std_logic;
  signal clk3c: std_logic;
  signal clk3d: std_logic;
  signal clk3e: std_logic;
  signal clk3f: std_logic;
  signal clk4a: std_logic;
  signal clk4b: std_logic;
  signal clk4c: std_logic;
  signal clk4d: std_logic;
  signal clk4e: std_logic;
  signal clk4f: std_logic;
  signal clk5: std_logic;
  signal clk5a: std_logic;
  signal dc0: std_logic;
  signal dc1: std_logic;
  signal dc2: std_logic;
  signal dc3: std_logic;
  signal dc4: std_logic;
  signal dc5: std_logic;
  signal dc6: std_logic;
  signal dc7: std_logic;
  signal dc8: std_logic;
  signal dc9: std_logic;
  signal dest: std_logic;
  signal destm: std_logic;
  signal destmd: std_logic;
  signal destspcd: std_logic;
  signal dispenb: std_logic;
  signal dn: std_logic;
  signal dp: std_logic;
  signal dparok: std_logic;
  signal dpc0: std_logic;
  signal dpc10: std_logic;
  signal dpc11: std_logic;
  signal dpc12: std_logic;
  signal dpc13: std_logic;
  signal dpc1: std_logic;
  signal dpc2: std_logic;
  signal dpc3: std_logic;
  signal dpc4: std_logic;
  signal dpc5: std_logic;
  signal dpc6: std_logic;
  signal dpc7: std_logic;
  signal dpc8: std_logic;
  signal dpc9: std_logic;
  signal dr: std_logic;
  signal err: std_logic;
  signal hi10: std_logic;
  signal hi11: std_logic;
  signal hi12: std_logic;
  signal hi1: std_logic;
  signal hi2: std_logic;
  signal hi3: std_logic;
  signal hi4: std_logic;
  signal hi5: std_logic;
  signal hi6: std_logic;
  signal hi7: std_logic;
  signal hi8: std_logic;
  signal hi9: std_logic;
  signal i0: std_logic;
  signal i10: std_logic;
  signal i11: std_logic;
  signal i12: std_logic;
  signal i13: std_logic;
  signal i14: std_logic;
  signal i15: std_logic;
  signal i16: std_logic;
  signal i17: std_logic;
  signal i18: std_logic;
  signal i19: std_logic;
  signal i1: std_logic;
  signal i20: std_logic;
  signal i21: std_logic;
  signal i22: std_logic;
  signal i23: std_logic;
  signal i24: std_logic;
  signal i25: std_logic;
  signal i26: std_logic;
  signal i27: std_logic;
  signal i28: std_logic;
  signal i29: std_logic;
  signal i2: std_logic;
  signal i30: std_logic;
  signal i31: std_logic;
  signal i32: std_logic;
  signal i33: std_logic;
  signal i34: std_logic;
  signal i35: std_logic;
  signal i36: std_logic;
  signal i37: std_logic;
  signal i38: std_logic;
  signal i39: std_logic;
  signal i3: std_logic;
  signal i40: std_logic;
  signal i41: std_logic;
  signal i42: std_logic;
  signal i43: std_logic;
  signal i44: std_logic;
  signal i45: std_logic;
  signal i46: std_logic;
  signal i47: std_logic;
  signal i48: std_logic;
  signal i4: std_logic;
  signal i5: std_logic;
  signal i6: std_logic;
  signal i7: std_logic;
  signal i8: std_logic;
  signal i9: std_logic;
  signal idebug: std_logic;
  signal imod: std_logic;
  signal imodd: std_logic;
  signal iparok: std_logic;
  signal ipc0: std_logic;
  signal ipc10: std_logic;
  signal ipc11: std_logic;
  signal ipc12: std_logic;
  signal ipc13: std_logic;
  signal ipc1: std_logic;
  signal ipc2: std_logic;
  signal ipc3: std_logic;
  signal ipc4: std_logic;
  signal ipc5: std_logic;
  signal ipc6: std_logic;
  signal ipc7: std_logic;
  signal ipc8: std_logic;
  signal ipc9: std_logic;
  signal ir0: std_logic;
  signal ir10: std_logic;
  signal ir11: std_logic;
  signal ir12: std_logic;
  signal ir13: std_logic;
  signal ir14: std_logic;
  signal ir15: std_logic;
  signal ir16: std_logic;
  signal ir17: std_logic;
  signal ir18: std_logic;
  signal ir19: std_logic;
  signal ir1: std_logic;
  signal ir20: std_logic;
  signal ir21: std_logic;
  signal ir22: std_logic;
  signal ir23: std_logic;
  signal ir24: std_logic;
  signal ir25: std_logic;
  signal ir26: std_logic;
  signal ir27: std_logic;
  signal ir28: std_logic;
  signal ir29: std_logic;
  signal ir2: std_logic;
  signal ir30: std_logic;
  signal ir31: std_logic;
  signal ir32: std_logic;
  signal ir33: std_logic;
  signal ir34: std_logic;
  signal ir35: std_logic;
  signal ir36: std_logic;
  signal ir37: std_logic;
  signal ir38: std_logic;
  signal ir39: std_logic;
  signal ir3: std_logic;
  signal ir40: std_logic;
  signal ir41: std_logic;
  signal ir42: std_logic;
  signal ir43: std_logic;
  signal ir44: std_logic;
  signal ir45: std_logic;
  signal ir46: std_logic;
  signal ir47: std_logic;
  signal ir48: std_logic;
  signal ir4: std_logic;
  signal ir5: std_logic;
  signal ir6: std_logic;
  signal ir7: std_logic;
  signal ir8: std_logic;
  signal ir9: std_logic;
  signal irdisp: std_logic;
  signal irjump: std_logic;
  signal iwr0: std_logic;
  signal iwr10: std_logic;
  signal iwr11: std_logic;
  signal iwr12: std_logic;
  signal iwr13: std_logic;
  signal iwr14: std_logic;
  signal iwr15: std_logic;
  signal iwr16: std_logic;
  signal iwr17: std_logic;
  signal iwr18: std_logic;
  signal iwr19: std_logic;
  signal iwr1: std_logic;
  signal iwr20: std_logic;
  signal iwr21: std_logic;
  signal iwr22: std_logic;
  signal iwr23: std_logic;
  signal iwr24: std_logic;
  signal iwr25: std_logic;
  signal iwr26: std_logic;
  signal iwr27: std_logic;
  signal iwr28: std_logic;
  signal iwr29: std_logic;
  signal iwr2: std_logic;
  signal iwr30: std_logic;
  signal iwr31: std_logic;
  signal iwr32: std_logic;
  signal iwr33: std_logic;
  signal iwr34: std_logic;
  signal iwr35: std_logic;
  signal iwr36: std_logic;
  signal iwr37: std_logic;
  signal iwr38: std_logic;
  signal iwr39: std_logic;
  signal iwr3: std_logic;
  signal iwr40: std_logic;
  signal iwr41: std_logic;
  signal iwr42: std_logic;
  signal iwr43: std_logic;
  signal iwr44: std_logic;
  signal iwr45: std_logic;
  signal iwr46: std_logic;
  signal iwr47: std_logic;
  signal iwr48: std_logic;
  signal iwr4: std_logic;
  signal iwr5: std_logic;
  signal iwr6: std_logic;
  signal iwr7: std_logic;
  signal iwr8: std_logic;
  signal iwr9: std_logic;
  signal iwrited: std_logic;
  signal jcond: std_logic;
  signal l0: std_logic;
  signal l10: std_logic;
  signal l11: std_logic;
  signal l12: std_logic;
  signal l13: std_logic;
  signal l14: std_logic;
  signal l15: std_logic;
  signal l16: std_logic;
  signal l17: std_logic;
  signal l18: std_logic;
  signal l19: std_logic;
  signal l1: std_logic;
  signal l20: std_logic;
  signal l21: std_logic;
  signal l22: std_logic;
  signal l23: std_logic;
  signal l24: std_logic;
  signal l25: std_logic;
  signal l26: std_logic;
  signal l27: std_logic;
  signal l28: std_logic;
  signal l29: std_logic;
  signal l2: std_logic;
  signal l30: std_logic;
  signal l31: std_logic;
  signal l3: std_logic;
  signal l4: std_logic;
  signal l5: std_logic;
  signal l6: std_logic;
  signal l7: std_logic;
  signal l8: std_logic;
  signal l9: std_logic;
  signal lc10: std_logic;
  signal lc11: std_logic;
  signal lc12: std_logic;
  signal lc13: std_logic;
  signal lc14: std_logic;
  signal lc15: std_logic;
  signal lc16: std_logic;
  signal lc17: std_logic;
  signal lc18: std_logic;
  signal lc19: std_logic;
  signal lc20: std_logic;
  signal lc21: std_logic;
  signal lc22: std_logic;
  signal lc23: std_logic;
  signal lc24: std_logic;
  signal lc25: std_logic;
  signal lc2: std_logic;
  signal lc3: std_logic;
  signal lc4: std_logic;
  signal lc5: std_logic;
  signal lc6: std_logic;
  signal lc7: std_logic;
  signal lc8: std_logic;
  signal lc9: std_logic;
  signal lcinc: std_logic;
  signal lcry3: std_logic;
  signal lparity: std_logic;
  signal m0: std_logic;
  signal m10: std_logic;
  signal m11: std_logic;
  signal m12: std_logic;
  signal m13: std_logic;
  signal m14: std_logic;
  signal m15: std_logic;
  signal m16: std_logic;
  signal m17: std_logic;
  signal m18: std_logic;
  signal m19: std_logic;
  signal m1: std_logic;
  signal m20: std_logic;
  signal m21: std_logic;
  signal m22: std_logic;
  signal m23: std_logic;
  signal m24: std_logic;
  signal m25: std_logic;
  signal m26: std_logic;
  signal m27: std_logic;
  signal m28: std_logic;
  signal m29: std_logic;
  signal m2: std_logic;
  signal m30: std_logic;
  signal m31: std_logic;
  signal m3: std_logic;
  signal m4: std_logic;
  signal m5: std_logic;
  signal m6: std_logic;
  signal m7: std_logic;
  signal m8: std_logic;
  signal m9: std_logic;
  signal machrun: std_logic;
  signal mapi10: std_logic;
  signal mapi11: std_logic;
  signal mapi12: std_logic;
  signal mapi13: std_logic;
  signal mapi14: std_logic;
  signal mapi15: std_logic;
  signal mapi16: std_logic;
  signal mapi17: std_logic;
  signal mapi18: std_logic;
  signal mapi19: std_logic;
  signal mapi20: std_logic;
  signal mapi21: std_logic;
  signal mapi22: std_logic;
  signal mapi23: std_logic;
  signal mapi8: std_logic;
  signal mapi9: std_logic;
  signal mclk1a: std_logic;
  signal mclk5: std_logic;
  signal mdhaspar: std_logic;
  signal mdpar: std_logic;
  signal mdparodd: std_logic;
  signal mdsela: std_logic;
  signal mdselb: std_logic;
  signal memparok: std_logic;
  signal memstart: std_logic;
  signal mf0: std_logic;
  signal mf10: std_logic;
  signal mf11: std_logic;
  signal mf12: std_logic;
  signal mf13: std_logic;
  signal mf14: std_logic;
  signal mf15: std_logic;
  signal mf16: std_logic;
  signal mf17: std_logic;
  signal mf18: std_logic;
  signal mf19: std_logic;
  signal mf1: std_logic;
  signal mf20: std_logic;
  signal mf21: std_logic;
  signal mf22: std_logic;
  signal mf23: std_logic;
  signal mf24: std_logic;
  signal mf25: std_logic;
  signal mf26: std_logic;
  signal mf27: std_logic;
  signal mf28: std_logic;
  signal mf29: std_logic;
  signal mf2: std_logic;
  signal mf30: std_logic;
  signal mf31: std_logic;
  signal mf3: std_logic;
  signal mf4: std_logic;
  signal mf5: std_logic;
  signal mf6: std_logic;
  signal mf7: std_logic;
  signal mf8: std_logic;
  signal mf9: std_logic;
  signal mmemparok: std_logic;
  signal mparity: std_logic;
  signal msk0: std_logic;
  signal msk10: std_logic;
  signal msk11: std_logic;
  signal msk12: std_logic;
  signal msk13: std_logic;
  signal msk14: std_logic;
  signal msk15: std_logic;
  signal msk16: std_logic;
  signal msk17: std_logic;
  signal msk18: std_logic;
  signal msk19: std_logic;
  signal msk1: std_logic;
  signal msk20: std_logic;
  signal msk21: std_logic;
  signal msk22: std_logic;
  signal msk23: std_logic;
  signal msk24: std_logic;
  signal msk25: std_logic;
  signal msk26: std_logic;
  signal msk27: std_logic;
  signal msk28: std_logic;
  signal msk29: std_logic;
  signal msk2: std_logic;
  signal msk30: std_logic;
  signal msk31: std_logic;
  signal msk3: std_logic;
  signal msk4: std_logic;
  signal msk5: std_logic;
  signal msk6: std_logic;
  signal msk7: std_logic;
  signal msk8: std_logic;
  signal msk9: std_logic;
  signal n: std_logic;
  signal needfetch: std_logic;
  signal nop: std_logic;
  signal ob0: std_logic;
  signal ob10: std_logic;
  signal ob11: std_logic;
  signal ob12: std_logic;
  signal ob13: std_logic;
  signal ob14: std_logic;
  signal ob15: std_logic;
  signal ob16: std_logic;
  signal ob17: std_logic;
  signal ob18: std_logic;
  signal ob19: std_logic;
  signal ob1: std_logic;
  signal ob20: std_logic;
  signal ob21: std_logic;
  signal ob22: std_logic;
  signal ob23: std_logic;
  signal ob24: std_logic;
  signal ob25: std_logic;
  signal ob26: std_logic;
  signal ob27: std_logic;
  signal ob28: std_logic;
  signal ob29: std_logic;
  signal ob2: std_logic;
  signal ob30: std_logic;
  signal ob31: std_logic;
  signal ob3: std_logic;
  signal ob4: std_logic;
  signal ob5: std_logic;
  signal ob6: std_logic;
  signal ob7: std_logic;
  signal ob8: std_logic;
  signal ob9: std_logic;
  signal opc0: std_logic;
  signal opc10: std_logic;
  signal opc11: std_logic;
  signal opc12: std_logic;
  signal opc13: std_logic;
  signal opc1: std_logic;
  signal opc2: std_logic;
  signal opc3: std_logic;
  signal opc4: std_logic;
  signal opc5: std_logic;
  signal opc6: std_logic;
  signal opc7: std_logic;
  signal opc8: std_logic;
  signal opc9: std_logic;
  signal opcclk: std_logic;
  signal osel0a: std_logic;
  signal osel0b: std_logic;
  signal osel1a: std_logic;
  signal osel1b: std_logic;
  signal pc0: std_logic;
  signal pc10: std_logic;
  signal pc11: std_logic;
  signal pc12: std_logic;
  signal pc13: std_logic;
  signal pc1: std_logic;
  signal pc2: std_logic;
  signal pc3: std_logic;
  signal pc4: std_logic;
  signal pc5: std_logic;
  signal pc6: std_logic;
  signal pc7: std_logic;
  signal pc8: std_logic;
  signal pc9: std_logic;
  signal pcs0: std_logic;
  signal pcs1: std_logic;
  signal pdlenb: std_logic;
  signal pdlparok: std_logic;
  signal pdlwrited: std_logic;
  signal promdisable: std_logic;
  signal promdisabled: std_logic;
  signal q0: std_logic;
  signal q31: std_logic;
  signal r0: std_logic;
  signal r10: std_logic;
  signal r11: std_logic;
  signal r12: std_logic;
  signal r13: std_logic;
  signal r14: std_logic;
  signal r15: std_logic;
  signal r16: std_logic;
  signal r17: std_logic;
  signal r18: std_logic;
  signal r19: std_logic;
  signal r1: std_logic;
  signal r20: std_logic;
  signal r21: std_logic;
  signal r22: std_logic;
  signal r23: std_logic;
  signal r24: std_logic;
  signal r25: std_logic;
  signal r26: std_logic;
  signal r27: std_logic;
  signal r28: std_logic;
  signal r29: std_logic;
  signal r2: std_logic;
  signal r30: std_logic;
  signal r31: std_logic;
  signal r3: std_logic;
  signal r4: std_logic;
  signal r5: std_logic;
  signal r6: std_logic;
  signal r7: std_logic;
  signal r8: std_logic;
  signal r9: std_logic;
  signal reset: std_logic;
  signal sintr: std_logic;
  signal spc0: std_logic;
  signal spc10: std_logic;
  signal spc11: std_logic;
  signal spc12: std_logic;
  signal spc13: std_logic;
  signal spc14: std_logic;
  signal spc1: std_logic;
  signal spc1a: std_logic;
  signal spc2: std_logic;
  signal spc3: std_logic;
  signal spc4: std_logic;
  signal spc5: std_logic;
  signal spc6: std_logic;
  signal spc7: std_logic;
  signal spc8: std_logic;
  signal spc9: std_logic;
  signal spcdrive: std_logic;
  signal spcenb: std_logic;
  signal spcparok: std_logic;
  signal spcwpass: std_logic;
  signal spush: std_logic;
  signal spushd: std_logic;
  signal spy0: std_logic;
  signal spy10: std_logic;
  signal spy11: std_logic;
  signal spy12: std_logic;
  signal spy13: std_logic;
  signal spy14: std_logic;
  signal spy15: std_logic;
  signal spy1: std_logic;
  signal spy2: std_logic;
  signal spy3: std_logic;
  signal spy4: std_logic;
  signal spy5: std_logic;
  signal spy6: std_logic;
  signal spy7: std_logic;
  signal spy8: std_logic;
  signal spy9: std_logic;
  signal srcm: std_logic;
  signal srcpdlidx: std_logic;
  signal srcpdlptr: std_logic;
  signal srun: std_logic;
  signal ssdone: std_logic;
  signal sspeed0: std_logic;
  signal sspeed1: std_logic;
  signal trapa: std_logic;
  signal trapb: std_logic;
  signal trapenb: std_logic;
  signal tse1a: std_logic;
  signal tse1b: std_logic;
  signal tse2: std_logic;
  signal tse3a: std_logic;
  signal tse4a: std_logic;
  signal tse4b: std_logic;
  signal v0parok: std_logic;
  signal vmasela: std_logic;
  signal vmaselb: std_logic;
  signal vmoparok: std_logic;
  signal wadr0: std_logic;
  signal wadr1: std_logic;
  signal wadr2: std_logic;
  signal wadr3: std_logic;
  signal wadr4: std_logic;
  signal wmapd: std_logic;
  signal wp1a: std_logic;
  signal wp1b: std_logic;
  signal wp2: std_logic;
  signal wp3a: std_logic;
  signal wp4a: std_logic;
  signal wp4b: std_logic;
  signal wp4c: std_logic;
begin
  alu_set_inst: alu_set port map (
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    a31b => a31b,
    \-div\ => \-div\,
    hi12 => hi12,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    \-ir12\ => \-ir12\,
    \-ir13\ => \-ir13\,
    \-iralu\ => \-iralu\,
    irjump => irjump,
    \-irjump\ => \-irjump\,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    \-mul\ => \-mul\,
    q0 => q0,
    a12 => a12,
    \a=m\ => \a=m\,
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    alu31 => alu31,
    alu32 => alu32,
    \-ir0\ => \-ir0\,
    \-ir1\ => \-ir1\,
    \-ir2\ => \-ir2\,
    \-ir3\ => \-ir3\,
    \-ir4\ => \-ir4\,
    osel0a => osel0a,
    osel0b => osel0b,
    osel1a => osel1a,
    osel1b => osel1b
  );
  amem_set_inst: amem_set port map (
    clk3d => clk3d,
    clk3e => clk3e,
    dest => dest,
    destm => destm,
    hi3 => hi3,
    hi5 => hi5,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
    \-reset\ => \-reset\,
    tse3a => tse3a,
    tse4a => tse4a,
    wp3a => wp3a,
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    a31b => a31b,
    aparity => aparity,
    destmd => destmd,
    wadr0 => wadr0,
    wadr1 => wadr1,
    wadr2 => wadr2,
    wadr3 => wadr3,
    wadr4 => wadr4
  );
  ampar_set_inst: ampar_set port map (
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31b => a31b,
    aparity => aparity,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    mparity => mparity,
    pdlenb => pdlenb,
    srcm => srcm,
    aparok => aparok,
    mmemparok => mmemparok,
    pdlparok => pdlparok
  );
  clock_set_inst: clock_set port map (
    \-clock reset b\ => \-clock reset b\,
    \-hang\ => \-hang\,
    hi1 => hi1,
    hi2 => hi2,
    hi3 => hi3,
    hi4 => hi4,
    hi5 => hi5,
    hi6 => hi6,
    hi7 => hi7,
    hi8 => hi8,
    hi9 => hi9,
    hi10 => hi10,
    hi11 => hi11,
    hi12 => hi12,
    \-ilong\ => \-ilong\,
    lcry3 => lcry3,
    machrun => machrun,
    \-machruna\ => \-machruna\,
    reset => reset,
    \-srcpdlidx\ => \-srcpdlidx\,
    \-srcpdlptr\ => \-srcpdlptr\,
    sspeed0 => sspeed0,
    sspeed1 => sspeed1,
    clk5 => clk5,
    clk1a => clk1a,
    clk2a => clk2a,
    clk2b => clk2b,
    clk2c => clk2c,
    clk3a => clk3a,
    clk3b => clk3b,
    clk3c => clk3c,
    clk3d => clk3d,
    clk3e => clk3e,
    clk3f => clk3f,
    clk4a => clk4a,
    clk4b => clk4b,
    clk4c => clk4c,
    clk4d => clk4d,
    clk4e => clk4e,
    clk4f => clk4f,
    \-clk2c\ => \-clk2c\,
    \-clk3g\ => \-clk3g\,
    \-clk4e\ => \-clk4e\,
    \-lcry3\ => \-lcry3\,
    mclk5 => mclk5,
    mclk1a => mclk1a,
    \-reset\ => \-reset\,
    srcpdlidx => srcpdlidx,
    srcpdlptr => srcpdlptr,
    \-tpr60\ => \-tpr60\,
    tse2 => tse2,
    tse1a => tse1a,
    tse1b => tse1b,
    tse3a => tse3a,
    tse4a => tse4a,
    tse4b => tse4b,
    \-upperhighok\ => \-upperhighok\,
    wp2 => wp2,
    wp1a => wp1a,
    wp1b => wp1b,
    wp3a => wp3a,
    wp4a => wp4a,
    wp4b => wp4b,
    wp4c => wp4c,
    \-wp5\ => \-wp5\
  );
  decode_set_inst: decode_set port map (
    hi5 => hi5,
    \-idebug\ => \-idebug\,
    ir3 => ir3,
    ir4 => ir4,
    ir8 => ir8,
    ir10 => ir10,
    ir11 => ir11,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir43 => ir43,
    ir44 => ir44,
    \-ir31\ => \-ir31\,
    nop => nop,
    dest => dest,
    \-destimod0\ => \-destimod0\,
    \-destimod1\ => \-destimod1\,
    \-destintctl\ => \-destintctl\,
    \-destlc\ => \-destlc\,
    destm => destm,
    \-destmdr\ => \-destmdr\,
    \-destmem\ => \-destmem\,
    \-destpdl(p)\ => \-destpdl(p)\,
    \-destpdl(x)\ => \-destpdl(x)\,
    \-destpdlp\ => \-destpdlp\,
    \-destpdltop\ => \-destpdltop\,
    \-destpdlx\ => \-destpdlx\,
    \-destspc\ => \-destspc\,
    \-destvma\ => \-destvma\,
    \-div\ => \-div\,
    \-funct2\ => \-funct2\,
    imod => imod,
    \-iralu\ => \-iralu\,
    \-irbyte\ => \-irbyte\,
    irdisp => irdisp,
    \-irdisp\ => \-irdisp\,
    irjump => irjump,
    \-irjump\ => \-irjump\,
    \-mul\ => \-mul\,
    \-srcdc\ => \-srcdc\,
    \-srclc\ => \-srclc\,
    \-srcmap\ => \-srcmap\,
    \-srcmd\ => \-srcmd\,
    \-srcopc\ => \-srcopc\,
    \-srcpdlidx\ => \-srcpdlidx\,
    \-srcpdlpop\ => \-srcpdlpop\,
    \-srcpdlptr\ => \-srcpdlptr\,
    \-srcpdltop\ => \-srcpdltop\,
    \-srcq\ => \-srcq\,
    \-srcspc\ => \-srcspc\,
    \-srcspcpop\ => \-srcspcpop\,
    \-srcvma\ => \-srcvma\
  );
  dmem_set_inst: dmem_set port map (
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    clk3e => clk3e,
    dispenb => dispenb,
    \-funct2\ => \-funct2\,
    hi4 => hi4,
    hi6 => hi6,
    hi11 => hi11,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    \-irdisp\ => \-irdisp\,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    wp2 => wp2,
    dn => dn,
    dpc0 => dpc0,
    dpc1 => dpc1,
    dpc2 => dpc2,
    dpc3 => dpc3,
    dpc5 => dpc5,
    dpc6 => dpc6,
    dpc7 => dpc7,
    dpc8 => dpc8,
    dpc9 => dpc9,
    dpc10 => dpc10,
    dpc11 => dpc11,
    dpc12 => dpc12,
    dpc13 => dpc13,
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    dc0 => dc0,
    dc1 => dc1,
    dc2 => dc2,
    dc3 => dc3,
    dc4 => dc4,
    dc5 => dc5,
    dc6 => dc6,
    dc7 => dc7,
    dc8 => dc8,
    dc9 => dc9,
    dp => dp,
    dparok => dparok,
    dpc4 => dpc4,
    dr => dr,
    \-vmo18\ => \-vmo18\,
    \-vmo19\ => \-vmo19\
  );
  fetch_set_inst: fetch_set port map (
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    clk2c => clk2c,
    clk4c => clk4c,
    \-idebug\ => \-idebug\,
    \-lddbirh\ => \-lddbirh\,
    \-lddbirl\ => \-lddbirl\,
    \-lddbirm\ => \-lddbirm\,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15,
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48
  );
  flowc_set_inst: flowc_set port map (
    clk3c => clk3c,
    dp => dp,
    dr => dr,
    \-funct2\ => \-funct2\,
    hi4 => hi4,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir42 => ir42,
    irdisp => irdisp,
    \-irdisp\ => \-irdisp\,
    irjump => irjump,
    jcond => jcond,
    \-jcond\ => \-jcond\,
    \-nop11\ => \-nop11\,
    \-reset\ => \-reset\,
    \-srcspc\ => \-srcspc\,
    \-srcspcpop\ => \-srcspcpop\,
    \-trap\ => \-trap\,
    tse3a => tse3a,
    wp4c => wp4c,
    \-destspc\ => \-destspc\,
    destspcd => destspcd,
    dispenb => dispenb,
    dn => dn,
    iwrited => iwrited,
    \-iwrited\ => \-iwrited\,
    n => n,
    nop => nop,
    \-nopa\ => \-nopa\,
    pcs0 => pcs0,
    pcs1 => pcs1,
    spcdrive => spcdrive,
    \-spcdrive\ => \-spcdrive\,
    spcenb => spcenb,
    \-spcnt\ => \-spcnt\,
    \-spcpass\ => \-spcpass\,
    spcwpass => spcwpass,
    \-spcwpass\ => \-spcwpass\,
    \-spop\ => \-spop\,
    spush => spush,
    spushd => spushd,
    \-srcspcpopreal\ => \-srcspcpopreal\,
    \-swpa\ => \-swpa\,
    \-swpb\ => \-swpb\
  );
  imem_set_inst: imem_set port map (
    hi1 => hi1,
    idebug => idebug,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    iwr32 => iwr32,
    iwr33 => iwr33,
    iwr34 => iwr34,
    iwr35 => iwr35,
    iwr36 => iwr36,
    iwr37 => iwr37,
    iwr38 => iwr38,
    iwr39 => iwr39,
    iwr40 => iwr40,
    iwr41 => iwr41,
    iwr42 => iwr42,
    iwr43 => iwr43,
    iwr44 => iwr44,
    iwr45 => iwr45,
    iwr46 => iwr46,
    iwr47 => iwr47,
    iwr48 => iwr48,
    \-iwrited\ => \-iwrited\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    promdisabled => promdisabled,
    \-wp5\ => \-wp5\,
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    \-iwriteda\ => \-iwriteda\,
    \-promdisabled\ => \-promdisabled\
  );
  ireg_set_inst: ireg_set port map (
    clk3a => clk3a,
    clk3b => clk3b,
    \-destimod0\ => \-destimod0\,
    \-destimod1\ => \-destimod1\,
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48,
    imodd => imodd,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    iparok => iparok,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir10 => ir10,
    ir11 => ir11,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    ir31 => ir31,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    ir42 => ir42,
    ir43 => ir43,
    ir44 => ir44,
    ir45 => ir45,
    ir46 => ir46,
    ir47 => ir47,
    ir48 => ir48
  );
  jumpc_set_inst: jumpc_set port map (
    \a=m\ => \a=m\,
    alu32 => alu32,
    clk3c => clk3c,
    \-destintctl\ => \-destintctl\,
    hi4 => hi4,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir5 => ir5,
    ir45 => ir45,
    ir46 => ir46,
    \-nopa\ => \-nopa\,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    r0 => r0,
    \-reset\ => \-reset\,
    sintr => sintr,
    \-vmaok\ => \-vmaok\,
    \-ilong\ => \-ilong\,
    \int.enable\ => \int.enable\,
    jcond => jcond,
    \-jcond\ => \-jcond\,
    \lc byte mode\ => \lc byte mode\,
    \prog.unibus.reset\ => \prog.unibus.reset\,
    \sequence.break\ => \sequence.break\,
    \-statbit\ => \-statbit\
  );
  lcreg_set_inst: lcreg_set port map (
    clk1a => clk1a,
    clk2a => clk2a,
    clk2c => clk2c,
    clk3c => clk3c,
    \-destlc\ => \-destlc\,
    hi11 => hi11,
    \int.enable\ => \int.enable\,
    ir10 => ir10,
    ir11 => ir11,
    ir24 => ir24,
    \-ir3\ => \-ir3\,
    \-ir4\ => \-ir4\,
    irdisp => irdisp,
    \lc byte mode\ => \lc byte mode\,
    \-lcry3\ => \-lcry3\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    \prog.unibus.reset\ => \prog.unibus.reset\,
    \-reset\ => \-reset\,
    \sequence.break\ => \sequence.break\,
    spc1 => spc1,
    spc14 => spc14,
    \-spop\ => \-spop\,
    \-srclc\ => \-srclc\,
    \-srcspcpopreal\ => \-srcspcpopreal\,
    tse1a => tse1a,
    \-ifetch\ => \-ifetch\,
    lc2 => lc2,
    lc3 => lc3,
    lc4 => lc4,
    lc5 => lc5,
    lc6 => lc6,
    lc7 => lc7,
    lc8 => lc8,
    lc9 => lc9,
    lc10 => lc10,
    lc11 => lc11,
    lc12 => lc12,
    lc13 => lc13,
    lc14 => lc14,
    lc15 => lc15,
    lc16 => lc16,
    lc17 => lc17,
    lc18 => lc18,
    lc19 => lc19,
    lc20 => lc20,
    lc21 => lc21,
    lc22 => lc22,
    lc23 => lc23,
    lc24 => lc24,
    lc25 => lc25,
    lcinc => lcinc,
    lcry3 => lcry3,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    needfetch => needfetch,
    \-sh3\ => \-sh3\,
    \-sh4\ => \-sh4\,
    sintr => sintr,
    spc1a => spc1a
  );
  lreg_set_inst: lreg_set port map (
    clk3f => clk3f,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity
  );
  md_set_inst: md_set port map (
    \-clk2c\ => \-clk2c\,
    \-destmdr\ => \-destmdr\,
    hi11 => hi11,
    mdparodd => mdparodd,
    mdsela => mdsela,
    mdselb => mdselb,
    \-memdrive.a\ => \-memdrive.a\,
    \-memdrive.b\ => \-memdrive.b\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    \-srcmd\ => \-srcmd\,
    tse2 => tse2,
    \-md0\ => \-md0\,
    \-md1\ => \-md1\,
    \-md2\ => \-md2\,
    \-md3\ => \-md3\,
    \-md4\ => \-md4\,
    \-md5\ => \-md5\,
    \-md6\ => \-md6\,
    \-md7\ => \-md7\,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-md24\ => \-md24\,
    \-md25\ => \-md25\,
    \-md26\ => \-md26\,
    \-md27\ => \-md27\,
    \-md28\ => \-md28\,
    \-md29\ => \-md29\,
    \-md30\ => \-md30\,
    \-md31\ => \-md31\,
    mdhaspar => mdhaspar,
    mdpar => mdpar,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31
  );
  mmem_set_inst: mmem_set port map (
    clk4a => clk4a,
    clk4e => clk4e,
    destmd => destmd,
    hi2 => hi2,
    hi3 => hi3,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    \-ir31\ => \-ir31\,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
    pdlenb => pdlenb,
    spcenb => spcenb,
    tse1a => tse1a,
    tse4a => tse4a,
    wadr0 => wadr0,
    wadr1 => wadr1,
    wadr2 => wadr2,
    wadr3 => wadr3,
    wadr4 => wadr4,
    wp4b => wp4b,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    mparity => mparity,
    srcm => srcm
  );
  mos_set_inst: mos_set port map (
    a0 => a0,
    a1 => a1,
    a2 => a2,
    a3 => a3,
    a4 => a4,
    a5 => a5,
    a6 => a6,
    a7 => a7,
    a8 => a8,
    a9 => a9,
    a10 => a10,
    a11 => a11,
    a12 => a12,
    a13 => a13,
    a14 => a14,
    a15 => a15,
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31b => a31b,
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    alu31 => alu31,
    alu32 => alu32,
    msk0 => msk0,
    msk1 => msk1,
    msk2 => msk2,
    msk3 => msk3,
    msk4 => msk4,
    msk5 => msk5,
    msk6 => msk6,
    msk7 => msk7,
    msk8 => msk8,
    msk9 => msk9,
    msk10 => msk10,
    msk11 => msk11,
    msk12 => msk12,
    msk13 => msk13,
    msk14 => msk14,
    msk15 => msk15,
    msk16 => msk16,
    msk17 => msk17,
    msk18 => msk18,
    msk19 => msk19,
    msk20 => msk20,
    msk21 => msk21,
    msk22 => msk22,
    msk23 => msk23,
    msk24 => msk24,
    msk25 => msk25,
    msk26 => msk26,
    msk27 => msk27,
    msk28 => msk28,
    msk29 => msk29,
    msk30 => msk30,
    msk31 => msk31,
    osel0a => osel0a,
    osel0b => osel0b,
    osel1a => osel1a,
    osel1b => osel1b,
    q31 => q31,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    r7 => r7,
    r8 => r8,
    r9 => r9,
    r10 => r10,
    r11 => r11,
    r12 => r12,
    r13 => r13,
    r14 => r14,
    r15 => r15,
    r16 => r16,
    r17 => r17,
    r18 => r18,
    r19 => r19,
    r20 => r20,
    r21 => r21,
    r22 => r22,
    r23 => r23,
    r24 => r24,
    r25 => r25,
    r26 => r26,
    r27 => r27,
    r28 => r28,
    r29 => r29,
    r30 => r30,
    r31 => r31,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31
  );
  npc_set_inst: npc_set port map (
    clk4b => clk4b,
    dpc4 => dpc4,
    hi4 => hi4,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    pcs0 => pcs0,
    pcs1 => pcs1,
    spc1a => spc1a,
    trapa => trapa,
    trapb => trapb,
    dpc0 => dpc0,
    dpc1 => dpc1,
    dpc2 => dpc2,
    dpc3 => dpc3,
    dpc5 => dpc5,
    dpc6 => dpc6,
    dpc7 => dpc7,
    dpc8 => dpc8,
    dpc9 => dpc9,
    dpc10 => dpc10,
    dpc11 => dpc11,
    dpc12 => dpc12,
    dpc13 => dpc13,
    ipc0 => ipc0,
    ipc1 => ipc1,
    ipc2 => ipc2,
    ipc3 => ipc3,
    ipc4 => ipc4,
    ipc5 => ipc5,
    ipc6 => ipc6,
    ipc7 => ipc7,
    ipc8 => ipc8,
    ipc9 => ipc9,
    ipc10 => ipc10,
    ipc11 => ipc11,
    ipc12 => ipc12,
    ipc13 => ipc13,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    spc0 => spc0,
    spc2 => spc2,
    spc3 => spc3,
    spc4 => spc4,
    spc5 => spc5,
    spc6 => spc6,
    spc7 => spc7,
    spc8 => spc8,
    spc9 => spc9,
    spc10 => spc10,
    spc11 => spc11,
    spc12 => spc12,
    spc13 => spc13
  );
  olord_set_inst: olord_set port map (
    aparok => aparok,
    clk5 => clk5,
    dparok => dparok,
    iparok => iparok,
    \-ldclk\ => \-ldclk\,
    \-ldopc\ => \-ldopc\,
    mclk5 => mclk5,
    memparok => memparok,
    mmemparok => mmemparok,
    pdlparok => pdlparok,
    spcparok => spcparok,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    \-stc32\ => \-stc32\,
    \-tpr60\ => \-tpr60\,
    \-upperhighok\ => \-upperhighok\,
    v0parok => v0parok,
    vmoparok => vmoparok,
    \-wait\ => \-wait\,
    \-ldmode\ => \-ldmode\,
    \-reset\ => \-reset\,
    \-ape\ => \-ape\,
    \boot.trap\ => \boot.trap\,
    \-clk5\ => \-clk5\,
    clk5a => clk5a,
    \-clock reset b\ => \-clock reset b\,
    \-dpe\ => \-dpe\,
    err => err,
    hi1 => hi1,
    hi2 => hi2,
    \-higherr\ => \-higherr\,
    idebug => idebug,
    \-idebug\ => \-idebug\,
    \-ipe\ => \-ipe\,
    \-ldstat\ => \-ldstat\,
    \lpc.hold\ => \lpc.hold\,
    machrun => machrun,
    \-machruna\ => \-machruna\,
    \-mempe\ => \-mempe\,
    \-mpe\ => \-mpe\,
    \-nop11\ => \-nop11\,
    opcclk => opcclk,
    \-opcinh\ => \-opcinh\,
    \-pdlpe\ => \-pdlpe\,
    promdisable => promdisable,
    promdisabled => promdisabled,
    reset => reset,
    \-spe\ => \-spe\,
    srun => srun,
    ssdone => ssdone,
    sspeed0 => sspeed0,
    sspeed1 => sspeed1,
    \-stathalt\ => \-stathalt\,
    trapenb => trapenb,
    \-v0pe\ => \-v0pe\,
    \-v1pe\ => \-v1pe\
  );
  opc_set_inst: opc_set port map (
    \-clk5\ => \-clk5\,
    dc0 => dc0,
    dc1 => dc1,
    dc2 => dc2,
    dc3 => dc3,
    dc4 => dc4,
    dc5 => dc5,
    dc6 => dc6,
    dc7 => dc7,
    dc8 => dc8,
    dc9 => dc9,
    hi2 => hi2,
    opcclk => opcclk,
    \-opcinh\ => \-opcinh\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    \-srcdc\ => \-srcdc\,
    \-srcopc\ => \-srcopc\,
    \-srcpdlidx\ => \-srcpdlidx\,
    \-srcpdlptr\ => \-srcpdlptr\,
    tse1b => tse1b,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    opc0 => opc0,
    opc1 => opc1,
    opc2 => opc2,
    opc3 => opc3,
    opc4 => opc4,
    opc5 => opc5,
    opc6 => opc6,
    opc7 => opc7,
    opc8 => opc8,
    opc9 => opc9,
    opc10 => opc10,
    opc11 => opc11,
    opc12 => opc12,
    opc13 => opc13
  );
  pdl_set_inst: pdl_set port map (
    clk3f => clk3f,
    clk4a => clk4a,
    clk4b => clk4b,
    clk4f => clk4f,
    \-clk4e\ => \-clk4e\,
    \-destpdl(p)\ => \-destpdl(p)\,
    \-destpdl(x)\ => \-destpdl(x)\,
    \-destpdlp\ => \-destpdlp\,
    \-destpdltop\ => \-destpdltop\,
    \-destpdlx\ => \-destpdlx\,
    \-destspc\ => \-destspc\,
    imod => imod,
    ir30 => ir30,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    l19 => l19,
    l20 => l20,
    l21 => l21,
    l22 => l22,
    l23 => l23,
    l24 => l24,
    l25 => l25,
    l26 => l26,
    l27 => l27,
    l28 => l28,
    l29 => l29,
    l30 => l30,
    l31 => l31,
    lparity => lparity,
    nop => nop,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    \-reset\ => \-reset\,
    srcpdlidx => srcpdlidx,
    \-srcpdlpop\ => \-srcpdlpop\,
    srcpdlptr => srcpdlptr,
    \-srcpdltop\ => \-srcpdltop\,
    tse4b => tse4b,
    wp4a => wp4a,
    imodd => imodd,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mparity => mparity,
    pdlenb => pdlenb,
    pdlwrited => pdlwrited
  );
  prom_set_inst: prom_set port map (
    \-ape\ => \-ape\,
    \-dpe\ => \-dpe\,
    hi2 => hi2,
    \-idebug\ => \-idebug\,
    \-ipe\ => \-ipe\,
    \-iwriteda\ => \-iwriteda\,
    \-mempe\ => \-mempe\,
    \-mpe\ => \-mpe\,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    \-pdlpe\ => \-pdlpe\,
    \-promdisabled\ => \-promdisabled\,
    \-spe\ => \-spe\,
    \-v0pe\ => \-v0pe\,
    \-v1pe\ => \-v1pe\,
    i0 => i0,
    i1 => i1,
    i2 => i2,
    i3 => i3,
    i4 => i4,
    i5 => i5,
    i6 => i6,
    i7 => i7,
    i8 => i8,
    i9 => i9,
    i10 => i10,
    i11 => i11,
    i12 => i12,
    i13 => i13,
    i14 => i14,
    i15 => i15,
    i16 => i16,
    i17 => i17,
    i18 => i18,
    i19 => i19,
    i20 => i20,
    i21 => i21,
    i22 => i22,
    i23 => i23,
    i24 => i24,
    i25 => i25,
    i26 => i26,
    i27 => i27,
    i28 => i28,
    i29 => i29,
    i30 => i30,
    i31 => i31,
    i32 => i32,
    i33 => i33,
    i34 => i34,
    i35 => i35,
    i36 => i36,
    i37 => i37,
    i38 => i38,
    i39 => i39,
    i40 => i40,
    i41 => i41,
    i42 => i42,
    i43 => i43,
    i44 => i44,
    i45 => i45,
    i46 => i46,
    i47 => i47,
    i48 => i48
  );
  qreg_set_inst: qreg_set port map (
    alu0 => alu0,
    alu1 => alu1,
    alu2 => alu2,
    alu3 => alu3,
    alu4 => alu4,
    alu5 => alu5,
    alu6 => alu6,
    alu7 => alu7,
    alu8 => alu8,
    alu9 => alu9,
    alu10 => alu10,
    alu11 => alu11,
    alu12 => alu12,
    alu13 => alu13,
    alu14 => alu14,
    alu15 => alu15,
    alu16 => alu16,
    alu17 => alu17,
    alu18 => alu18,
    alu19 => alu19,
    alu20 => alu20,
    alu21 => alu21,
    alu22 => alu22,
    alu23 => alu23,
    alu24 => alu24,
    alu25 => alu25,
    alu26 => alu26,
    alu27 => alu27,
    alu28 => alu28,
    alu29 => alu29,
    alu30 => alu30,
    alu31 => alu31,
    clk2b => clk2b,
    hi7 => hi7,
    \-ir0\ => \-ir0\,
    \-ir1\ => \-ir1\,
    \-iralu\ => \-iralu\,
    \-srcq\ => \-srcq\,
    tse2 => tse2,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    q0 => q0,
    q31 => q31
  );
  shifter_masker_set_inst: shifter_masker_set port map (
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    \-ir0\ => \-ir0\,
    ir12 => ir12,
    ir13 => ir13,
    \-ir1\ => \-ir1\,
    \-ir2\ => \-ir2\,
    ir31 => ir31,
    \-irbyte\ => \-irbyte\,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    \-sh3\ => \-sh3\,
    \-sh4\ => \-sh4\,
    \a=m\ => \a=m\,
    \-ir12\ => \-ir12\,
    \-ir13\ => \-ir13\,
    \-ir31\ => \-ir31\,
    m5 => m5,
    msk0 => msk0,
    msk1 => msk1,
    msk2 => msk2,
    msk3 => msk3,
    msk4 => msk4,
    msk5 => msk5,
    msk6 => msk6,
    msk7 => msk7,
    msk8 => msk8,
    msk9 => msk9,
    msk10 => msk10,
    msk11 => msk11,
    msk12 => msk12,
    msk13 => msk13,
    msk14 => msk14,
    msk15 => msk15,
    msk16 => msk16,
    msk17 => msk17,
    msk18 => msk18,
    msk19 => msk19,
    msk20 => msk20,
    msk21 => msk21,
    msk22 => msk22,
    msk23 => msk23,
    msk24 => msk24,
    msk25 => msk25,
    msk26 => msk26,
    msk27 => msk27,
    msk28 => msk28,
    msk29 => msk29,
    msk30 => msk30,
    msk31 => msk31,
    r0 => r0,
    r1 => r1,
    r2 => r2,
    r3 => r3,
    r4 => r4,
    r5 => r5,
    r6 => r6,
    r7 => r7,
    r8 => r8,
    r9 => r9,
    r10 => r10,
    r11 => r11,
    r12 => r12,
    r13 => r13,
    r14 => r14,
    r15 => r15,
    r16 => r16,
    r17 => r17,
    r18 => r18,
    r19 => r19,
    r20 => r20,
    r21 => r21,
    r22 => r22,
    r23 => r23,
    r24 => r24,
    r25 => r25,
    r26 => r26,
    r27 => r27,
    r28 => r28,
    r29 => r29,
    r30 => r30,
    r31 => r31
  );
  spc_set_inst: spc_set port map (
    clk4b => clk4b,
    clk4c => clk4c,
    clk4d => clk4d,
    clk4f => clk4f,
    destspcd => destspcd,
    ipc0 => ipc0,
    ipc1 => ipc1,
    ipc2 => ipc2,
    ipc3 => ipc3,
    ipc4 => ipc4,
    ipc5 => ipc5,
    ipc6 => ipc6,
    ipc7 => ipc7,
    ipc8 => ipc8,
    ipc9 => ipc9,
    ipc10 => ipc10,
    ipc11 => ipc11,
    ipc12 => ipc12,
    ipc13 => ipc13,
    ir25 => ir25,
    irdisp => irdisp,
    l0 => l0,
    l1 => l1,
    l2 => l2,
    l3 => l3,
    l4 => l4,
    l5 => l5,
    l6 => l6,
    l7 => l7,
    l8 => l8,
    l9 => l9,
    l10 => l10,
    l11 => l11,
    l12 => l12,
    l13 => l13,
    l14 => l14,
    l15 => l15,
    l16 => l16,
    l17 => l17,
    l18 => l18,
    \lpc.hold\ => \lpc.hold\,
    n => n,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    spcdrive => spcdrive,
    \-spcdrive\ => \-spcdrive\,
    \-spcnt\ => \-spcnt\,
    \-spcpass\ => \-spcpass\,
    spcwpass => spcwpass,
    \-spcwpass\ => \-spcwpass\,
    spush => spush,
    \-swpa\ => \-swpa\,
    \-swpb\ => \-swpb\,
    hi1 => hi1,
    spc0 => spc0,
    spc2 => spc2,
    spc3 => spc3,
    spc4 => spc4,
    spc5 => spc5,
    spc6 => spc6,
    spc7 => spc7,
    spc8 => spc8,
    spc9 => spc9,
    spc10 => spc10,
    spc11 => spc11,
    spc12 => spc12,
    spc13 => spc13,
    hi2 => hi2,
    hi3 => hi3,
    hi4 => hi4,
    hi5 => hi5,
    hi6 => hi6,
    hi7 => hi7,
    hi8 => hi8,
    hi9 => hi9,
    hi10 => hi10,
    hi11 => hi11,
    hi12 => hi12,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    spc1 => spc1,
    spc14 => spc14,
    spcparok => spcparok
  );
  spy_set_inst: spy_set port map (
    a16 => a16,
    a17 => a17,
    a18 => a18,
    a19 => a19,
    a20 => a20,
    a21 => a21,
    a22 => a22,
    a23 => a23,
    a24 => a24,
    a25 => a25,
    a26 => a26,
    a27 => a27,
    a28 => a28,
    a29 => a29,
    a30 => a30,
    a31a => a31a,
    aa0 => aa0,
    aa1 => aa1,
    aa2 => aa2,
    aa3 => aa3,
    aa4 => aa4,
    aa5 => aa5,
    aa6 => aa6,
    aa7 => aa7,
    aa8 => aa8,
    aa9 => aa9,
    aa10 => aa10,
    aa11 => aa11,
    aa12 => aa12,
    aa13 => aa13,
    aa14 => aa14,
    aa15 => aa15,
    \-ape\ => \-ape\,
    destspcd => destspcd,
    \-dpe\ => \-dpe\,
    err => err,
    hi1 => hi1,
    \-higherr\ => \-higherr\,
    imodd => imodd,
    \-ipe\ => \-ipe\,
    ir0 => ir0,
    ir1 => ir1,
    ir2 => ir2,
    ir3 => ir3,
    ir4 => ir4,
    ir5 => ir5,
    ir6 => ir6,
    ir7 => ir7,
    ir8 => ir8,
    ir9 => ir9,
    ir10 => ir10,
    ir11 => ir11,
    ir12 => ir12,
    ir13 => ir13,
    ir14 => ir14,
    ir15 => ir15,
    ir16 => ir16,
    ir17 => ir17,
    ir18 => ir18,
    ir19 => ir19,
    ir20 => ir20,
    ir21 => ir21,
    ir22 => ir22,
    ir23 => ir23,
    ir24 => ir24,
    ir25 => ir25,
    ir26 => ir26,
    ir27 => ir27,
    ir28 => ir28,
    ir29 => ir29,
    ir30 => ir30,
    ir31 => ir31,
    ir32 => ir32,
    ir33 => ir33,
    ir34 => ir34,
    ir35 => ir35,
    ir36 => ir36,
    ir37 => ir37,
    ir38 => ir38,
    ir39 => ir39,
    ir40 => ir40,
    ir41 => ir41,
    ir42 => ir42,
    ir43 => ir43,
    ir44 => ir44,
    ir45 => ir45,
    ir46 => ir46,
    ir47 => ir47,
    ir48 => ir48,
    iwrited => iwrited,
    jcond => jcond,
    m0 => m0,
    m1 => m1,
    m2 => m2,
    m3 => m3,
    m4 => m4,
    m5 => m5,
    m6 => m6,
    m7 => m7,
    m8 => m8,
    m9 => m9,
    m10 => m10,
    m11 => m11,
    m12 => m12,
    m13 => m13,
    m14 => m14,
    m15 => m15,
    m16 => m16,
    m17 => m17,
    m18 => m18,
    m19 => m19,
    m20 => m20,
    m21 => m21,
    m22 => m22,
    m23 => m23,
    m24 => m24,
    m25 => m25,
    m26 => m26,
    m27 => m27,
    m28 => m28,
    m29 => m29,
    m30 => m30,
    m31 => m31,
    \-mempe\ => \-mempe\,
    \-mpe\ => \-mpe\,
    nop => nop,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    opc0 => opc0,
    opc1 => opc1,
    opc2 => opc2,
    opc3 => opc3,
    opc4 => opc4,
    opc5 => opc5,
    opc6 => opc6,
    opc7 => opc7,
    opc8 => opc8,
    opc9 => opc9,
    opc10 => opc10,
    opc11 => opc11,
    opc12 => opc12,
    opc13 => opc13,
    pc0 => pc0,
    pc1 => pc1,
    pc2 => pc2,
    pc3 => pc3,
    pc4 => pc4,
    pc5 => pc5,
    pc6 => pc6,
    pc7 => pc7,
    pc8 => pc8,
    pc9 => pc9,
    pc10 => pc10,
    pc11 => pc11,
    pc12 => pc12,
    pc13 => pc13,
    pcs0 => pcs0,
    pcs1 => pcs1,
    \-pdlpe\ => \-pdlpe\,
    pdlwrited => pdlwrited,
    promdisable => promdisable,
    \-spe\ => \-spe\,
    spushd => spushd,
    srun => srun,
    ssdone => ssdone,
    \-stathalt\ => \-stathalt\,
    \-v0pe\ => \-v0pe\,
    \-v1pe\ => \-v1pe\,
    \-vmaok\ => \-vmaok\,
    \-wait\ => \-wait\,
    wmapd => wmapd,
    \-ldclk\ => \-ldclk\,
    \-lddbirh\ => \-lddbirh\,
    \-lddbirl\ => \-lddbirl\,
    \-lddbirm\ => \-lddbirm\,
    \-ldmode\ => \-ldmode\,
    \-ldopc\ => \-ldopc\,
    \-spy.sth\ => \-spy.sth\,
    \-spy.stl\ => \-spy.stl\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15
  );
  stat_set_inst: stat_set port map (
    clk5a => clk5a,
    hi1 => hi1,
    iwr0 => iwr0,
    iwr1 => iwr1,
    iwr2 => iwr2,
    iwr3 => iwr3,
    iwr4 => iwr4,
    iwr5 => iwr5,
    iwr6 => iwr6,
    iwr7 => iwr7,
    iwr8 => iwr8,
    iwr9 => iwr9,
    iwr10 => iwr10,
    iwr11 => iwr11,
    iwr12 => iwr12,
    iwr13 => iwr13,
    iwr14 => iwr14,
    iwr15 => iwr15,
    iwr16 => iwr16,
    iwr17 => iwr17,
    iwr18 => iwr18,
    iwr19 => iwr19,
    iwr20 => iwr20,
    iwr21 => iwr21,
    iwr22 => iwr22,
    iwr23 => iwr23,
    iwr24 => iwr24,
    iwr25 => iwr25,
    iwr26 => iwr26,
    iwr27 => iwr27,
    iwr28 => iwr28,
    iwr29 => iwr29,
    iwr30 => iwr30,
    iwr31 => iwr31,
    \-ldstat\ => \-ldstat\,
    \-spy.sth\ => \-spy.sth\,
    \-spy.stl\ => \-spy.stl\,
    \-statbit\ => \-statbit\,
    spy0 => spy0,
    spy1 => spy1,
    spy2 => spy2,
    spy3 => spy3,
    spy4 => spy4,
    spy5 => spy5,
    spy6 => spy6,
    spy7 => spy7,
    spy8 => spy8,
    spy9 => spy9,
    spy10 => spy10,
    spy11 => spy11,
    spy12 => spy12,
    spy13 => spy13,
    spy14 => spy14,
    spy15 => spy15,
    \-stc32\ => \-stc32\
  );
  trap_set_inst: trap_set port map (
    \boot.trap\ => \boot.trap\,
    \-md0\ => \-md0\,
    \-md1\ => \-md1\,
    \-md2\ => \-md2\,
    \-md3\ => \-md3\,
    \-md4\ => \-md4\,
    \-md5\ => \-md5\,
    \-md6\ => \-md6\,
    \-md7\ => \-md7\,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-md24\ => \-md24\,
    \-md25\ => \-md25\,
    \-md26\ => \-md26\,
    \-md27\ => \-md27\,
    \-md28\ => \-md28\,
    \-md29\ => \-md29\,
    \-md30\ => \-md30\,
    \-md31\ => \-md31\,
    mdhaspar => mdhaspar,
    mdpar => mdpar,
    trapenb => trapenb,
    \use.md\ => \use.md\,
    \-wait\ => \-wait\,
    mdparodd => mdparodd,
    memparok => memparok,
    \-trap\ => \-trap\,
    trapa => trapa,
    trapb => trapb
  );
  vctl_set_inst: vctl_set port map (
    clk2a => clk2a,
    clk2c => clk2c,
    \-clk3g\ => \-clk3g\,
    \-destmdr\ => \-destmdr\,
    \-destmem\ => \-destmem\,
    \-destvma\ => \-destvma\,
    hi4 => hi4,
    hi11 => hi11,
    \-ifetch\ => \-ifetch\,
    ir19 => ir19,
    ir20 => ir20,
    lcinc => lcinc,
    \-lvmo22\ => \-lvmo22\,
    \-lvmo23\ => \-lvmo23\,
    mclk1a => mclk1a,
    needfetch => needfetch,
    \-nopa\ => \-nopa\,
    \-reset\ => \-reset\,
    \-srcmd\ => \-srcmd\,
    \-vma25\ => \-vma25\,
    \-vma26\ => \-vma26\,
    wp1a => wp1a,
    wp1b => wp1b,
    \-hang\ => \-hang\,
    mdsela => mdsela,
    mdselb => mdselb,
    \-memdrive.a\ => \-memdrive.a\,
    \-memdrive.b\ => \-memdrive.b\,
    memstart => memstart,
    \-memstart\ => \-memstart\,
    \-pfr\ => \-pfr\,
    \-pfw\ => \-pfw\,
    \use.md\ => \use.md\,
    \-vm0wpa\ => \-vm0wpa\,
    \-vm0wpb\ => \-vm0wpb\,
    \-vm1wpa\ => \-vm1wpa\,
    \-vm1wpb\ => \-vm1wpb\,
    \-vmaenb\ => \-vmaenb\,
    \-vmaok\ => \-vmaok\,
    vmasela => vmasela,
    vmaselb => vmaselb,
    \-wait\ => \-wait\,
    wmapd => wmapd
  );
  vma_set_inst: vma_set port map (
    clk1a => clk1a,
    clk2a => clk2a,
    clk2c => clk2c,
    lc2 => lc2,
    lc3 => lc3,
    lc4 => lc4,
    lc5 => lc5,
    lc6 => lc6,
    lc7 => lc7,
    lc8 => lc8,
    lc9 => lc9,
    lc10 => lc10,
    lc11 => lc11,
    lc12 => lc12,
    lc13 => lc13,
    lc14 => lc14,
    lc15 => lc15,
    lc16 => lc16,
    lc17 => lc17,
    lc18 => lc18,
    lc19 => lc19,
    lc20 => lc20,
    lc21 => lc21,
    lc22 => lc22,
    lc23 => lc23,
    lc24 => lc24,
    lc25 => lc25,
    \-md8\ => \-md8\,
    \-md9\ => \-md9\,
    \-md10\ => \-md10\,
    \-md11\ => \-md11\,
    \-md12\ => \-md12\,
    \-md13\ => \-md13\,
    \-md14\ => \-md14\,
    \-md15\ => \-md15\,
    \-md16\ => \-md16\,
    \-md17\ => \-md17\,
    \-md18\ => \-md18\,
    \-md19\ => \-md19\,
    \-md20\ => \-md20\,
    \-md21\ => \-md21\,
    \-md22\ => \-md22\,
    \-md23\ => \-md23\,
    \-memstart\ => \-memstart\,
    ob0 => ob0,
    ob1 => ob1,
    ob2 => ob2,
    ob3 => ob3,
    ob4 => ob4,
    ob5 => ob5,
    ob6 => ob6,
    ob7 => ob7,
    ob8 => ob8,
    ob9 => ob9,
    ob10 => ob10,
    ob11 => ob11,
    ob12 => ob12,
    ob13 => ob13,
    ob14 => ob14,
    ob15 => ob15,
    ob16 => ob16,
    ob17 => ob17,
    ob18 => ob18,
    ob19 => ob19,
    ob20 => ob20,
    ob21 => ob21,
    ob22 => ob22,
    ob23 => ob23,
    ob24 => ob24,
    ob25 => ob25,
    ob26 => ob26,
    ob27 => ob27,
    ob28 => ob28,
    ob29 => ob29,
    ob30 => ob30,
    ob31 => ob31,
    \-srcvma\ => \-srcvma\,
    tse2 => tse2,
    \-vmaenb\ => \-vmaenb\,
    vmasela => vmasela,
    vmaselb => vmaselb,
    mapi8 => mapi8,
    mapi9 => mapi9,
    mapi10 => mapi10,
    mapi11 => mapi11,
    mapi12 => mapi12,
    mapi13 => mapi13,
    mapi14 => mapi14,
    mapi15 => mapi15,
    mapi16 => mapi16,
    mapi17 => mapi17,
    mapi18 => mapi18,
    mapi19 => mapi19,
    mapi20 => mapi20,
    mapi21 => mapi21,
    mapi22 => mapi22,
    mapi23 => mapi23,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    \-vma0\ => \-vma0\,
    \-vma1\ => \-vma1\,
    \-vma2\ => \-vma2\,
    \-vma3\ => \-vma3\,
    \-vma4\ => \-vma4\,
    \-vma5\ => \-vma5\,
    \-vma6\ => \-vma6\,
    \-vma7\ => \-vma7\,
    \-vma8\ => \-vma8\,
    \-vma9\ => \-vma9\,
    \-vma10\ => \-vma10\,
    \-vma11\ => \-vma11\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    \-vma25\ => \-vma25\,
    \-vma26\ => \-vma26\,
    \-vma27\ => \-vma27\,
    \-vma28\ => \-vma28\,
    \-vma29\ => \-vma29\,
    \-vma30\ => \-vma30\,
    \-vma31\ => \-vma31\
  );
  vmaps_set_inst: vmaps_set port map (
    hi12 => hi12,
    mapi8 => mapi8,
    mapi9 => mapi9,
    mapi10 => mapi10,
    mapi11 => mapi11,
    mapi12 => mapi12,
    mapi13 => mapi13,
    mapi14 => mapi14,
    mapi15 => mapi15,
    mapi16 => mapi16,
    mapi17 => mapi17,
    mapi18 => mapi18,
    mapi19 => mapi19,
    mapi20 => mapi20,
    mapi21 => mapi21,
    mapi22 => mapi22,
    mapi23 => mapi23,
    memstart => memstart,
    \-pfr\ => \-pfr\,
    \-pfw\ => \-pfw\,
    \-srcmap\ => \-srcmap\,
    tse1a => tse1a,
    \-vm0wpa\ => \-vm0wpa\,
    \-vm0wpb\ => \-vm0wpb\,
    \-vm1wpa\ => \-vm1wpa\,
    \-vm1wpb\ => \-vm1wpb\,
    \-vma0\ => \-vma0\,
    \-vma1\ => \-vma1\,
    \-vma2\ => \-vma2\,
    \-vma3\ => \-vma3\,
    \-vma4\ => \-vma4\,
    \-vma5\ => \-vma5\,
    \-vma6\ => \-vma6\,
    \-vma7\ => \-vma7\,
    \-vma8\ => \-vma8\,
    \-vma9\ => \-vma9\,
    \-vma10\ => \-vma10\,
    \-vma11\ => \-vma11\,
    \-vma12\ => \-vma12\,
    \-vma13\ => \-vma13\,
    \-vma14\ => \-vma14\,
    \-vma15\ => \-vma15\,
    \-vma16\ => \-vma16\,
    \-vma17\ => \-vma17\,
    \-vma18\ => \-vma18\,
    \-vma19\ => \-vma19\,
    \-vma20\ => \-vma20\,
    \-vma21\ => \-vma21\,
    \-vma22\ => \-vma22\,
    \-vma23\ => \-vma23\,
    \-vma27\ => \-vma27\,
    \-vma28\ => \-vma28\,
    \-vma29\ => \-vma29\,
    \-vma30\ => \-vma30\,
    \-vma31\ => \-vma31\,
    \-vmo18\ => \-vmo18\,
    \-vmo19\ => \-vmo19\,
    \-lvmo22\ => \-lvmo22\,
    \-lvmo23\ => \-lvmo23\,
    mf0 => mf0,
    mf1 => mf1,
    mf2 => mf2,
    mf3 => mf3,
    mf4 => mf4,
    mf5 => mf5,
    mf6 => mf6,
    mf7 => mf7,
    mf8 => mf8,
    mf9 => mf9,
    mf10 => mf10,
    mf11 => mf11,
    mf12 => mf12,
    mf13 => mf13,
    mf14 => mf14,
    mf15 => mf15,
    mf16 => mf16,
    mf17 => mf17,
    mf18 => mf18,
    mf19 => mf19,
    mf20 => mf20,
    mf21 => mf21,
    mf22 => mf22,
    mf23 => mf23,
    mf24 => mf24,
    mf25 => mf25,
    mf26 => mf26,
    mf27 => mf27,
    mf28 => mf28,
    mf29 => mf29,
    mf30 => mf30,
    mf31 => mf31,
    v0parok => v0parok,
    vmoparok => vmoparok
  );
end architecture;
