library ieee;
use ieee.std_logic_1164.all;

entity cadr_spclch is
  port (
    \-spcdrive\     : in     std_logic;
    \-spcpass\      : in     std_logic;
    \-spcwpass\     : in     std_logic;
    clk4c           : in     std_logic;
    clk4d           : in     std_logic;
    hi1             : in     std_logic;
    spcdrive        : in     std_logic;
    spco0           : in     std_logic;
    spco1           : in     std_logic;
    spco10          : in     std_logic;
    spco11          : in     std_logic;
    spco12          : in     std_logic;
    spco13          : in     std_logic;
    spco14          : in     std_logic;
    spco15          : in     std_logic;
    spco16          : in     std_logic;
    spco17          : in     std_logic;
    spco18          : in     std_logic;
    spco2           : in     std_logic;
    spco3           : in     std_logic;
    spco4           : in     std_logic;
    spco5           : in     std_logic;
    spco6           : in     std_logic;
    spco7           : in     std_logic;
    spco8           : in     std_logic;
    spco9           : in     std_logic;
    spcopar         : in     std_logic;
    spcptr0         : in     std_logic;
    spcptr1         : in     std_logic;
    spcptr2         : in     std_logic;
    spcptr3         : in     std_logic;
    spcptr4         : in     std_logic;
    spcw0           : in     std_logic;
    spcw1           : in     std_logic;
    spcw10          : in     std_logic;
    spcw11          : in     std_logic;
    spcw12          : in     std_logic;
    spcw13          : in     std_logic;
    spcw14          : in     std_logic;
    spcw15          : in     std_logic;
    spcw16          : in     std_logic;
    spcw17          : in     std_logic;
    spcw18          : in     std_logic;
    spcw2           : in     std_logic;
    spcw3           : in     std_logic;
    spcw4           : in     std_logic;
    spcw5           : in     std_logic;
    spcw6           : in     std_logic;
    spcw7           : in     std_logic;
    spcw8           : in     std_logic;
    spcw9           : in     std_logic;
    spcwpar         : in     std_logic;
    spcwpass        : in     std_logic;
    m0              : out    std_logic;
    m1              : out    std_logic;
    m10             : out    std_logic;
    m11             : out    std_logic;
    m12             : out    std_logic;
    m13             : out    std_logic;
    m14             : out    std_logic;
    m15             : out    std_logic;
    m16             : out    std_logic;
    m17             : out    std_logic;
    m18             : out    std_logic;
    m19             : out    std_logic;
    m2              : out    std_logic;
    m20             : out    std_logic;
    m21             : out    std_logic;
    m22             : out    std_logic;
    m23             : out    std_logic;
    m24             : out    std_logic;
    m25             : out    std_logic;
    m26             : out    std_logic;
    m27             : out    std_logic;
    m28             : out    std_logic;
    m29             : out    std_logic;
    m3              : out    std_logic;
    m30             : out    std_logic;
    m31             : out    std_logic;
    m4              : out    std_logic;
    m5              : out    std_logic;
    m6              : out    std_logic;
    m7              : out    std_logic;
    m8              : out    std_logic;
    m9              : out    std_logic;
    spc0            : out    std_logic;
    spc1            : out    std_logic;
    spc10           : out    std_logic;
    spc11           : out    std_logic;
    spc12           : out    std_logic;
    spc13           : out    std_logic;
    spc14           : out    std_logic;
    spc15           : out    std_logic;
    spc16           : out    std_logic;
    spc17           : out    std_logic;
    spc18           : out    std_logic;
    spc2            : out    std_logic;
    spc3            : out    std_logic;
    spc4            : out    std_logic;
    spc5            : out    std_logic;
    spc6            : out    std_logic;
    spc7            : out    std_logic;
    spc8            : out    std_logic;
    spc9            : out    std_logic;
    spcpar          : out    std_logic
  );
end entity;
