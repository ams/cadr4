library ieee;
use ieee.std_logic_1164.all;

entity cadr_iram01 is
  port (
    pc0b     : out std_logic;
    pc1b     : out std_logic;
    pc2b     : out std_logic;
    pc3b     : out std_logic;
    pc4b     : out std_logic;
    pc5b     : out std_logic;
    i10      : out std_logic;
    \-iweb\  : in  std_logic;
    \-ice1a\ : in  std_logic;
    iwr10    : in  std_logic;
    pc11b    : out std_logic;
    pc10b    : out std_logic;
    pc9b     : out std_logic;
    pc8b     : out std_logic;
    pc7b     : out std_logic;
    pc6b     : out std_logic;
    i11      : out std_logic;
    iwr11    : in  std_logic;
    \-pcb6\  : in  std_logic;
    \-pcb7\  : in  std_logic;
    \-pcb8\  : in  std_logic;
    \-pcb9\  : in  std_logic;
    \-pcb10\ : in  std_logic;
    \-pcb11\ : in  std_logic;
    \-pcb0\  : in  std_logic;
    \-pcb1\  : in  std_logic;
    \-pcb2\  : in  std_logic;
    \-pcb3\  : in  std_logic;
    \-pcb4\  : in  std_logic;
    \-pcb5\  : in  std_logic;
    i5       : out std_logic;
    iwr5     : in  std_logic;
    i6       : out std_logic;
    iwr6     : in  std_logic;
    i7       : out std_logic;
    iwr7     : in  std_logic;
    i8       : out std_logic;
    iwr8     : in  std_logic;
    i9       : out std_logic;
    iwr9     : in  std_logic;
    i0       : out std_logic;
    iwr0     : in  std_logic;
    i1       : out std_logic;
    iwr1     : in  std_logic;
    i2       : out std_logic;
    iwr2     : in  std_logic;
    i3       : out std_logic;
    iwr3     : in  std_logic;
    i4       : out std_logic;
    iwr4     : in  std_logic);
end;
