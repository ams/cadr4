library ieee;
use ieee.std_logic_1164.all;

entity cadr_alatch is
  port (
    \-amemenb\      : in     std_logic;
    \-apassenb\     : in     std_logic;
    amem0           : in     std_logic;
    amem1           : in     std_logic;
    amem10          : in     std_logic;
    amem11          : in     std_logic;
    amem12          : in     std_logic;
    amem13          : in     std_logic;
    amem14          : in     std_logic;
    amem15          : in     std_logic;
    amem16          : in     std_logic;
    amem17          : in     std_logic;
    amem18          : in     std_logic;
    amem19          : in     std_logic;
    amem2           : in     std_logic;
    amem20          : in     std_logic;
    amem21          : in     std_logic;
    amem22          : in     std_logic;
    amem23          : in     std_logic;
    amem24          : in     std_logic;
    amem25          : in     std_logic;
    amem26          : in     std_logic;
    amem27          : in     std_logic;
    amem28          : in     std_logic;
    amem29          : in     std_logic;
    amem3           : in     std_logic;
    amem30          : in     std_logic;
    amem31          : in     std_logic;
    amem4           : in     std_logic;
    amem5           : in     std_logic;
    amem6           : in     std_logic;
    amem7           : in     std_logic;
    amem8           : in     std_logic;
    amem9           : in     std_logic;
    amemparity      : in     std_logic;
    apassenb        : in     std_logic;
    clk3e           : in     std_logic;
    hi5             : in     std_logic;
    l0              : in     std_logic;
    l1              : in     std_logic;
    l10             : in     std_logic;
    l11             : in     std_logic;
    l12             : in     std_logic;
    l13             : in     std_logic;
    l14             : in     std_logic;
    l15             : in     std_logic;
    l16             : in     std_logic;
    l17             : in     std_logic;
    l18             : in     std_logic;
    l19             : in     std_logic;
    l2              : in     std_logic;
    l20             : in     std_logic;
    l21             : in     std_logic;
    l22             : in     std_logic;
    l23             : in     std_logic;
    l24             : in     std_logic;
    l25             : in     std_logic;
    l26             : in     std_logic;
    l27             : in     std_logic;
    l28             : in     std_logic;
    l29             : in     std_logic;
    l3              : in     std_logic;
    l30             : in     std_logic;
    l31             : in     std_logic;
    l4              : in     std_logic;
    l5              : in     std_logic;
    l6              : in     std_logic;
    l7              : in     std_logic;
    l8              : in     std_logic;
    l9              : in     std_logic;
    lparity         : in     std_logic;
    a0              : out    std_logic;
    a1              : out    std_logic;
    a10             : out    std_logic;
    a11             : out    std_logic;
    a12             : out    std_logic;
    a13             : out    std_logic;
    a14             : out    std_logic;
    a15             : out    std_logic;
    a16             : out    std_logic;
    a17             : out    std_logic;
    a18             : out    std_logic;
    a19             : out    std_logic;
    a2              : out    std_logic;
    a20             : out    std_logic;
    a21             : out    std_logic;
    a22             : out    std_logic;
    a23             : out    std_logic;
    a24             : out    std_logic;
    a25             : out    std_logic;
    a26             : out    std_logic;
    a27             : out    std_logic;
    a28             : out    std_logic;
    a29             : out    std_logic;
    a3              : out    std_logic;
    a30             : out    std_logic;
    a31a            : out    std_logic;
    a31b            : out    std_logic;
    a4              : out    std_logic;
    a5              : out    std_logic;
    a6              : out    std_logic;
    a7              : out    std_logic;
    a8              : out    std_logic;
    a9              : out    std_logic;
    aparity         : out    std_logic
  );
end entity cadr_alatch;
