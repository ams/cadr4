library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_spc is
  port (
    \-swpa\   : in  std_logic;
    gnd       : in  std_logic;
    spcw14    : in  std_logic;
    spcptr4   : out std_logic;
    hi1       : out std_logic;
    spco14    : out std_logic;
    spco15    : out std_logic;
    spcptr3   : out std_logic;
    spcptr2   : out std_logic;
    spcptr1   : out std_logic;
    spcptr0   : out std_logic;
    spcw15    : in  std_logic;
    spcw12    : in  std_logic;
    spco12    : out std_logic;
    spco13    : out std_logic;
    spcw13    : in  std_logic;
    spcw10    : in  std_logic;
    spco10    : out std_logic;
    spco11    : out std_logic;
    spcw11    : in  std_logic;
    spcopar   : out std_logic;
    spco18    : out std_logic;
    spco17    : out std_logic;
    spco16    : out std_logic;
    hi2       : out std_logic;
    hi3       : out std_logic;
    hi4       : out std_logic;
    hi5       : out std_logic;
    hi6       : out std_logic;
    hi7       : out std_logic;
    \-swpb\   : in  std_logic;
    spcw4     : in  std_logic;
    spco4     : out std_logic;
    spco5     : out std_logic;
    spcw5     : in  std_logic;
    spcw2     : in  std_logic;
    spco2     : out std_logic;
    spco3     : out std_logic;
    spcw3     : in  std_logic;
    spcw0     : in  std_logic;
    spco0     : out std_logic;
    spco1     : out std_logic;
    spcw1     : in  std_logic;
    spco9     : out std_logic;
    spco8     : out std_logic;
    spco7     : out std_logic;
    spco6     : out std_logic;
    hi8       : out std_logic;
    hi9       : out std_logic;
    hi10      : out std_logic;
    hi11      : out std_logic;
    hi12      : out std_logic;
    spush     : in  std_logic;
    clk4f     : in  std_logic;
    \-spcnt\  : in  std_logic;
    \-spccry\ : out std_logic;
    spcw18    : in  std_logic;
    spcwpar   : in  std_logic;
    spcw16    : in  std_logic;
    spcw17    : in  std_logic;
    spcw8     : in  std_logic;
    spcw9     : in  std_logic;
    spcw6     : in  std_logic;
    spcw7     : in  std_logic);
end;

architecture ttl of cadr_spc is
  signal nc182 : std_logic;
  signal nc183 : std_logic;
  signal nc184 : std_logic;
  signal nc185 : std_logic;
  signal nc186 : std_logic;
  signal nc187 : std_logic;
  signal nc188 : std_logic;
  signal nc189 : std_logic;
  signal nc190 : std_logic;
  signal nc191 : std_logic;
  signal nc192 : std_logic;
  signal nc193 : std_logic;
  signal nc194 : std_logic;
  signal nc195 : std_logic;
begin
  spc_4e21 : dm82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw14, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco14, d1 => spco15, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw15, we1_n => gnd);
  spc_4e22 : dm82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw12, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco12, d1 => spco13, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw13, we1_n => gnd);
  spc_4e23 : dm82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw10, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco10, d1 => spco11, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw11, we1_n => gnd);
  spc_4e24 : res20 port map(r2       => spcopar, r3 => spco18, r4 => spco17, r5 => spco16, r6 => spco15, r7 => hi1, r8 => hi2, r9 => hi3, r11 => hi4, r12 => hi5, r13 => hi6, r14 => hi7, r15 => spco14, r16 => spco13, r17 => spco12, r18 => spco11, r19 => spco10);
  spc_4e26 : dm82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw4, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco4, d1 => spco5, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw5, we1_n => gnd);
  spc_4e27 : dm82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw2, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco2, d1 => spco3, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw3, we1_n => gnd);
  spc_4e28 : dm82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw0, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco0, d1 => spco1, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw1, we1_n => gnd);
  spc_4e29 : res20 port map(r2       => spco9, r3 => spco8, r4 => spco7, r5 => spco6, r6 => spco5, r7 => hi8, r8 => hi9, r9 => hi10, r11 => hi11, r12 => hi12, r13 => nc182, r14 => nc183, r15 => spco4, r16 => spco3, r17 => spco2, r18 => spco1, r19 => spco0);
  spc_4f23 : sn74s169 port map(up_dn => spush, clk => clk4f, i0 => nc192, i1 => nc193, i2 => nc194, i3 => nc195, enb_p_n => gnd, load_n => hi1, enb_t_n => \-spcnt\, o3 => spcptr3, o2 => spcptr2, o1 => spcptr1, o0 => spcptr0, co_n => \-spccry\);
  spc_4f24 : dm82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw18, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco18, d1 => spcopar, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcwpar, we1_n => gnd);
  spc_4f25 : dm82s21 port map(wclk_n => \-swpa\, we0_n => gnd, i0 => spcw16, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco16, d1 => spco17, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw17, we1_n => gnd);
  spc_4f28 : sn74s169 port map(up_dn => spush, clk => clk4f, i0 => nc184, i1 => nc185, i2 => nc186, i3 => nc187, enb_p_n => gnd, load_n => hi1, enb_t_n => \-spccry\, o3 => nc188, o2 => nc189, o1 => nc190, o0 => spcptr4, co_n => nc191);
  spc_4f29 : dm82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw8, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco8, d1 => spco9, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw9, we1_n => gnd);
  spc_4f30 : dm82s21 port map(wclk_n => \-swpb\, we0_n => gnd, i0 => spcw6, a4 => spcptr4, ce => hi1, strobe => hi1, d0 => spco6, d1 => spco7, a3 => spcptr3, a2 => spcptr2, a1 => spcptr1, a0 => spcptr0, i1 => spcw7, we1_n => gnd);
end architecture;
