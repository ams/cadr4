library ieee;
use ieee.std_logic_1164.all;

library ttl;
use ttl.sn74.all;
use ttl.other.all;

library cadr;
use cadr.utilities.all;

entity cadr_shift0 is
  port (
    m5    : out std_logic;
    m6    : in  std_logic;
    m7    : in  std_logic;
    m8    : in  std_logic;
    m9    : in  std_logic;
    m10   : in  std_logic;
    m11   : in  std_logic;
    s1    : in  std_logic;
    s0    : in  std_logic;
    sa11  : out std_logic;
    sa10  : out std_logic;
    gnd   : in  std_logic;
    sa9   : out std_logic;
    sa8   : out std_logic;
    m29   : in  std_logic;
    m30   : in  std_logic;
    m31   : in  std_logic;
    m0    : in  std_logic;
    m1    : in  std_logic;
    m2    : in  std_logic;
    m3    : in  std_logic;
    sa3   : out std_logic;
    sa2   : out std_logic;
    sa1   : out std_logic;
    sa0   : out std_logic;
    m12   : in  std_logic;
    m13   : in  std_logic;
    m14   : in  std_logic;
    m15   : in  std_logic;
    sa15  : out std_logic;
    sa14  : out std_logic;
    sa13  : out std_logic;
    sa12  : out std_logic;
    m4    : in  std_logic;
    sa7   : out std_logic;
    sa6   : out std_logic;
    sa5   : out std_logic;
    sa4   : out std_logic;
    sa18  : in  std_logic;
    sa22  : in  std_logic;
    sa26  : in  std_logic;
    sa30  : in  std_logic;
    s3a   : in  std_logic;
    s2a   : in  std_logic;
    r14   : out std_logic;
    r10   : out std_logic;
    \-s4\ : in  std_logic;
    r6    : out std_logic;
    r2    : out std_logic;
    s4    : in  std_logic;
    sa19  : in  std_logic;
    sa23  : in  std_logic;
    sa27  : in  std_logic;
    sa31  : in  std_logic;
    r15   : out std_logic;
    r11   : out std_logic;
    r7    : out std_logic;
    r3    : out std_logic;
    sa16  : in  std_logic;
    sa20  : in  std_logic;
    sa24  : in  std_logic;
    sa28  : in  std_logic;
    r12   : out std_logic;
    r8    : out std_logic;
    r4    : out std_logic;
    r0    : out std_logic;
    sa17  : in  std_logic;
    sa21  : in  std_logic;
    sa25  : in  std_logic;
    sa29  : in  std_logic;
    r13   : out std_logic;
    r9    : out std_logic;
    r5    : out std_logic;
    r1    : out std_logic);
end;

architecture ttl of cadr_shift0 is
begin
  shift0_2c21 : am25s10 port map(i_3 => m5, i_2 => m6, i_1 => m7, i0 => m8, i1 => m9, i2 => m10, i3 => m11, sel1 => s1, sel0 => s0, o3 => sa11, o2 => sa10, ce_n => gnd, o1 => sa9, o0 => sa8);
  shift0_2c26 : am25s10 port map(i_3 => m29, i_2 => m30, i_1 => m31, i0 => m0, i1 => m1, i2 => m2, i3 => m3, sel1 => s1, sel0 => s0, o3 => sa3, o2 => sa2, ce_n => gnd, o1 => sa1, o0 => sa0);
  shift0_2d25 : am25s10 port map(i_3 => m9, i_2 => m10, i_1 => m11, i0 => m12, i1 => m13, i2 => m14, i3 => m15, sel1 => s1, sel0 => s0, o3 => sa15, o2 => sa14, ce_n => gnd, o1 => sa13, o0 => sa12);
  shift0_2d30 : am25s10 port map(i_3 => m1, i_2 => m2, i_1 => m3, i0 => m4, i1 => m5, i2 => m6, i3 => m7, sel1 => s1, sel0 => s0, o3 => sa7, o2 => sa6, ce_n => gnd, o1 => sa5, o0 => sa4);
  shift0_2e21 : am25s10 port map(i_3 => sa6, i_2 => sa10, i_1 => sa14, i0 => sa18, i1 => sa22, i2 => sa26, i3 => sa30, sel1 => s3a, sel0 => s2a, o3 => r14, o2 => r10, ce_n => \-s4\, o1 => r6, o0 => r2);
  shift0_2e22 : am25s10 port map(i_3 => sa22, i_2 => sa26, i_1 => sa30, i0 => sa2, i1 => sa6, i2 => sa10, i3 => sa14, sel1 => s3a, sel0 => s2a, o3 => r14, o2 => r10, ce_n => s4, o1 => r6, o0 => r2);
  shift0_2e23 : am25s10 port map(i_3 => sa7, i_2 => sa11, i_1 => sa15, i0 => sa19, i1 => sa23, i2 => sa27, i3 => sa31, sel1 => s3a, sel0 => s2a, o3 => r15, o2 => r11, ce_n => \-s4\, o1 => r7, o0 => r3);
  shift0_2e24 : am25s10 port map(i_3 => sa23, i_2 => sa27, i_1 => sa31, i0 => sa3, i1 => sa7, i2 => sa11, i3 => sa15, sel1 => s3a, sel0 => s2a, o3 => r15, o2 => r11, ce_n => s4, o1 => r7, o0 => r3);
  shift0_2e26 : am25s10 port map(i_3 => sa4, i_2 => sa8, i_1 => sa12, i0 => sa16, i1 => sa20, i2 => sa24, i3 => sa28, sel1 => s3a, sel0 => s2a, o3 => r12, o2 => r8, ce_n => \-s4\, o1 => r4, o0 => r0);
  shift0_2e27 : am25s10 port map(i_3 => sa20, i_2 => sa24, i_1 => sa28, i0 => sa0, i1 => sa4, i2 => sa8, i3 => sa12, sel1 => s3a, sel0 => s2a, o3 => r12, o2 => r8, ce_n => s4, o1 => r4, o0 => r0);
  shift0_2e28 : am25s10 port map(i_3 => sa5, i_2 => sa9, i_1 => sa13, i0 => sa17, i1 => sa21, i2 => sa25, i3 => sa29, sel1 => s3a, sel0 => s2a, o3 => r13, o2 => r9, ce_n => \-s4\, o1 => r5, o0 => r1);
  shift0_2e29 : am25s10 port map(i_3 => sa21, i_2 => sa25, i_1 => sa29, i0 => sa1, i1 => sa5, i2 => sa9, i3 => sa13, sel1 => s3a, sel0 => s2a, o3 => r13, o2 => r9, ce_n => s4, o1 => r5, o0 => r1);
end architecture;
