library ieee;
use ieee.std_logic_1164.all;

entity cadr_mo0 is
  port (
    a0              : in     std_logic;
    a1              : in     std_logic;
    a10             : in     std_logic;
    a11             : in     std_logic;
    a12             : in     std_logic;
    a13             : in     std_logic;
    a14             : in     std_logic;
    a15             : in     std_logic;
    a2              : in     std_logic;
    a3              : in     std_logic;
    a4              : in     std_logic;
    a5              : in     std_logic;
    a6              : in     std_logic;
    a7              : in     std_logic;
    a8              : in     std_logic;
    a9              : in     std_logic;
    alu0            : in     std_logic;
    alu1            : in     std_logic;
    alu10           : in     std_logic;
    alu11           : in     std_logic;
    alu12           : in     std_logic;
    alu13           : in     std_logic;
    alu14           : in     std_logic;
    alu15           : in     std_logic;
    alu16           : in     std_logic;
    alu2            : in     std_logic;
    alu3            : in     std_logic;
    alu4            : in     std_logic;
    alu5            : in     std_logic;
    alu6            : in     std_logic;
    alu7            : in     std_logic;
    alu8            : in     std_logic;
    alu9            : in     std_logic;
    msk0            : in     std_logic;
    msk1            : in     std_logic;
    msk10           : in     std_logic;
    msk11           : in     std_logic;
    msk12           : in     std_logic;
    msk13           : in     std_logic;
    msk14           : in     std_logic;
    msk15           : in     std_logic;
    msk2            : in     std_logic;
    msk3            : in     std_logic;
    msk4            : in     std_logic;
    msk5            : in     std_logic;
    msk6            : in     std_logic;
    msk7            : in     std_logic;
    msk8            : in     std_logic;
    msk9            : in     std_logic;
    osel0b          : in     std_logic;
    osel1b          : in     std_logic;
    q31             : in     std_logic;
    r0              : in     std_logic;
    r1              : in     std_logic;
    r10             : in     std_logic;
    r11             : in     std_logic;
    r12             : in     std_logic;
    r13             : in     std_logic;
    r14             : in     std_logic;
    r15             : in     std_logic;
    r2              : in     std_logic;
    r3              : in     std_logic;
    r4              : in     std_logic;
    r5              : in     std_logic;
    r6              : in     std_logic;
    r7              : in     std_logic;
    r8              : in     std_logic;
    r9              : in     std_logic;
    ob0             : out    std_logic;
    ob1             : out    std_logic;
    ob10            : out    std_logic;
    ob11            : out    std_logic;
    ob12            : out    std_logic;
    ob13            : out    std_logic;
    ob14            : out    std_logic;
    ob15            : out    std_logic;
    ob2             : out    std_logic;
    ob3             : out    std_logic;
    ob4             : out    std_logic;
    ob5             : out    std_logic;
    ob6             : out    std_logic;
    ob7             : out    std_logic;
    ob8             : out    std_logic;
    ob9             : out    std_logic
  );
end entity cadr_mo0;
