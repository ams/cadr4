library ieee;
use ieee.std_logic_1164.all;

entity spy4 is
  port (
    \-spy.flag1\ : out std_logic;
    \-wait\      : in  std_logic;
    spy8         : out std_logic;
    \-v1pe\      : in  std_logic;
    spy9         : out std_logic;
    \-v0pe\      : in  std_logic;
    spy10        : out std_logic;
    promdisable  : in  std_logic;
    spy11        : out std_logic;
    \-stathalt\  : in  std_logic;
    spy12        : out std_logic;
    err          : in  std_logic;
    spy13        : out std_logic;
    ssdone       : in  std_logic;
    spy14        : out std_logic;
    srun         : in  std_logic;
    spy15        : out std_logic;
    \-higherr\   : in  std_logic;
    spy0         : out std_logic;
    \-mempe\     : in  std_logic;
    spy1         : out std_logic;
    \-ipe\       : in  std_logic;
    spy2         : out std_logic;
    \-dpe\       : in  std_logic;
    spy3         : out std_logic;
    \-spe\       : in  std_logic;
    spy4         : out std_logic;
    \-pdlpe\     : in  std_logic;
    spy5         : out std_logic;
    \-mpe\       : in  std_logic;
    spy6         : out std_logic;
    \-ape\       : in  std_logic;
    spy7         : out std_logic;
    \-spy.pc\    : in  std_logic;
    gnd          : in  std_logic;
    pc13         : in  std_logic;
    pc12         : in  std_logic;
    pc11         : in  std_logic;
    pc10         : in  std_logic;
    pc9          : in  std_logic;
    pc8          : in  std_logic;
    pc7          : in  std_logic;
    pc6          : in  std_logic;
    pc5          : in  std_logic;
    pc4          : in  std_logic;
    pc3          : in  std_logic;
    pc2          : in  std_logic;
    pc1          : in  std_logic;
    pc0          : in  std_logic;
    \-spy.opc\   : in  std_logic;
    opc13        : in  std_logic;
    opc12        : in  std_logic;
    opc11        : in  std_logic;
    opc10        : in  std_logic;
    opc9         : in  std_logic;
    opc8         : in  std_logic;
    opc7         : in  std_logic;
    opc6         : in  std_logic;
    opc5         : in  std_logic;
    opc4         : in  std_logic;
    opc3         : in  std_logic;
    opc2         : in  std_logic;
    opc1         : in  std_logic;
    opc0         : in  std_logic);
end;
